magic
tech gf180mcuC
magscale 1 5
timestamp 1670151550
<< obsm1 >>
rect 672 855 149296 148273
<< metal2 >>
rect 2184 149600 2240 150000
rect 3472 149600 3528 150000
rect 4760 149600 4816 150000
rect 6048 149600 6104 150000
rect 7336 149600 7392 150000
rect 8624 149600 8680 150000
rect 9912 149600 9968 150000
rect 11200 149600 11256 150000
rect 12488 149600 12544 150000
rect 13776 149600 13832 150000
rect 15064 149600 15120 150000
rect 16352 149600 16408 150000
rect 17640 149600 17696 150000
rect 18928 149600 18984 150000
rect 20216 149600 20272 150000
rect 21504 149600 21560 150000
rect 22792 149600 22848 150000
rect 24080 149600 24136 150000
rect 25368 149600 25424 150000
rect 26656 149600 26712 150000
rect 27944 149600 28000 150000
rect 29232 149600 29288 150000
rect 30520 149600 30576 150000
rect 31808 149600 31864 150000
rect 33096 149600 33152 150000
rect 34384 149600 34440 150000
rect 35672 149600 35728 150000
rect 36960 149600 37016 150000
rect 38248 149600 38304 150000
rect 39536 149600 39592 150000
rect 40824 149600 40880 150000
rect 42112 149600 42168 150000
rect 43400 149600 43456 150000
rect 44688 149600 44744 150000
rect 45976 149600 46032 150000
rect 47264 149600 47320 150000
rect 48552 149600 48608 150000
rect 49840 149600 49896 150000
rect 51128 149600 51184 150000
rect 52416 149600 52472 150000
rect 53704 149600 53760 150000
rect 54992 149600 55048 150000
rect 56280 149600 56336 150000
rect 57568 149600 57624 150000
rect 58856 149600 58912 150000
rect 60144 149600 60200 150000
rect 61432 149600 61488 150000
rect 62720 149600 62776 150000
rect 64008 149600 64064 150000
rect 65296 149600 65352 150000
rect 66584 149600 66640 150000
rect 67872 149600 67928 150000
rect 69160 149600 69216 150000
rect 70448 149600 70504 150000
rect 71736 149600 71792 150000
rect 73024 149600 73080 150000
rect 74312 149600 74368 150000
rect 75600 149600 75656 150000
rect 76888 149600 76944 150000
rect 78176 149600 78232 150000
rect 79464 149600 79520 150000
rect 80752 149600 80808 150000
rect 82040 149600 82096 150000
rect 83328 149600 83384 150000
rect 84616 149600 84672 150000
rect 85904 149600 85960 150000
rect 87192 149600 87248 150000
rect 88480 149600 88536 150000
rect 89768 149600 89824 150000
rect 91056 149600 91112 150000
rect 92344 149600 92400 150000
rect 93632 149600 93688 150000
rect 94920 149600 94976 150000
rect 96208 149600 96264 150000
rect 97496 149600 97552 150000
rect 98784 149600 98840 150000
rect 100072 149600 100128 150000
rect 101360 149600 101416 150000
rect 102648 149600 102704 150000
rect 103936 149600 103992 150000
rect 105224 149600 105280 150000
rect 106512 149600 106568 150000
rect 107800 149600 107856 150000
rect 109088 149600 109144 150000
rect 110376 149600 110432 150000
rect 111664 149600 111720 150000
rect 112952 149600 113008 150000
rect 114240 149600 114296 150000
rect 115528 149600 115584 150000
rect 116816 149600 116872 150000
rect 118104 149600 118160 150000
rect 119392 149600 119448 150000
rect 120680 149600 120736 150000
rect 121968 149600 122024 150000
rect 123256 149600 123312 150000
rect 124544 149600 124600 150000
rect 125832 149600 125888 150000
rect 127120 149600 127176 150000
rect 128408 149600 128464 150000
rect 129696 149600 129752 150000
rect 130984 149600 131040 150000
rect 132272 149600 132328 150000
rect 133560 149600 133616 150000
rect 134848 149600 134904 150000
rect 136136 149600 136192 150000
rect 137424 149600 137480 150000
rect 138712 149600 138768 150000
rect 140000 149600 140056 150000
rect 141288 149600 141344 150000
rect 142576 149600 142632 150000
rect 143864 149600 143920 150000
rect 145152 149600 145208 150000
rect 146440 149600 146496 150000
rect 147728 149600 147784 150000
rect 6048 0 6104 400
rect 6328 0 6384 400
rect 6608 0 6664 400
rect 6888 0 6944 400
rect 7168 0 7224 400
rect 7448 0 7504 400
rect 7728 0 7784 400
rect 8008 0 8064 400
rect 8288 0 8344 400
rect 8568 0 8624 400
rect 8848 0 8904 400
rect 9128 0 9184 400
rect 9408 0 9464 400
rect 9688 0 9744 400
rect 9968 0 10024 400
rect 10248 0 10304 400
rect 10528 0 10584 400
rect 10808 0 10864 400
rect 11088 0 11144 400
rect 11368 0 11424 400
rect 11648 0 11704 400
rect 11928 0 11984 400
rect 12208 0 12264 400
rect 12488 0 12544 400
rect 12768 0 12824 400
rect 13048 0 13104 400
rect 13328 0 13384 400
rect 13608 0 13664 400
rect 13888 0 13944 400
rect 14168 0 14224 400
rect 14448 0 14504 400
rect 14728 0 14784 400
rect 15008 0 15064 400
rect 15288 0 15344 400
rect 15568 0 15624 400
rect 15848 0 15904 400
rect 16128 0 16184 400
rect 16408 0 16464 400
rect 16688 0 16744 400
rect 16968 0 17024 400
rect 17248 0 17304 400
rect 17528 0 17584 400
rect 17808 0 17864 400
rect 18088 0 18144 400
rect 18368 0 18424 400
rect 18648 0 18704 400
rect 18928 0 18984 400
rect 19208 0 19264 400
rect 19488 0 19544 400
rect 19768 0 19824 400
rect 20048 0 20104 400
rect 20328 0 20384 400
rect 20608 0 20664 400
rect 20888 0 20944 400
rect 21168 0 21224 400
rect 21448 0 21504 400
rect 21728 0 21784 400
rect 22008 0 22064 400
rect 22288 0 22344 400
rect 22568 0 22624 400
rect 22848 0 22904 400
rect 23128 0 23184 400
rect 23408 0 23464 400
rect 23688 0 23744 400
rect 23968 0 24024 400
rect 24248 0 24304 400
rect 24528 0 24584 400
rect 24808 0 24864 400
rect 25088 0 25144 400
rect 25368 0 25424 400
rect 25648 0 25704 400
rect 25928 0 25984 400
rect 26208 0 26264 400
rect 26488 0 26544 400
rect 26768 0 26824 400
rect 27048 0 27104 400
rect 27328 0 27384 400
rect 27608 0 27664 400
rect 27888 0 27944 400
rect 28168 0 28224 400
rect 28448 0 28504 400
rect 28728 0 28784 400
rect 29008 0 29064 400
rect 29288 0 29344 400
rect 29568 0 29624 400
rect 29848 0 29904 400
rect 30128 0 30184 400
rect 30408 0 30464 400
rect 30688 0 30744 400
rect 30968 0 31024 400
rect 31248 0 31304 400
rect 31528 0 31584 400
rect 31808 0 31864 400
rect 32088 0 32144 400
rect 32368 0 32424 400
rect 32648 0 32704 400
rect 32928 0 32984 400
rect 33208 0 33264 400
rect 33488 0 33544 400
rect 33768 0 33824 400
rect 34048 0 34104 400
rect 34328 0 34384 400
rect 34608 0 34664 400
rect 34888 0 34944 400
rect 35168 0 35224 400
rect 35448 0 35504 400
rect 35728 0 35784 400
rect 36008 0 36064 400
rect 36288 0 36344 400
rect 36568 0 36624 400
rect 36848 0 36904 400
rect 37128 0 37184 400
rect 37408 0 37464 400
rect 37688 0 37744 400
rect 37968 0 38024 400
rect 38248 0 38304 400
rect 38528 0 38584 400
rect 38808 0 38864 400
rect 39088 0 39144 400
rect 39368 0 39424 400
rect 39648 0 39704 400
rect 39928 0 39984 400
rect 40208 0 40264 400
rect 40488 0 40544 400
rect 40768 0 40824 400
rect 41048 0 41104 400
rect 41328 0 41384 400
rect 41608 0 41664 400
rect 41888 0 41944 400
rect 42168 0 42224 400
rect 42448 0 42504 400
rect 42728 0 42784 400
rect 43008 0 43064 400
rect 43288 0 43344 400
rect 43568 0 43624 400
rect 43848 0 43904 400
rect 44128 0 44184 400
rect 44408 0 44464 400
rect 44688 0 44744 400
rect 44968 0 45024 400
rect 45248 0 45304 400
rect 45528 0 45584 400
rect 45808 0 45864 400
rect 46088 0 46144 400
rect 46368 0 46424 400
rect 46648 0 46704 400
rect 46928 0 46984 400
rect 47208 0 47264 400
rect 47488 0 47544 400
rect 47768 0 47824 400
rect 48048 0 48104 400
rect 48328 0 48384 400
rect 48608 0 48664 400
rect 48888 0 48944 400
rect 49168 0 49224 400
rect 49448 0 49504 400
rect 49728 0 49784 400
rect 50008 0 50064 400
rect 50288 0 50344 400
rect 50568 0 50624 400
rect 50848 0 50904 400
rect 51128 0 51184 400
rect 51408 0 51464 400
rect 51688 0 51744 400
rect 51968 0 52024 400
rect 52248 0 52304 400
rect 52528 0 52584 400
rect 52808 0 52864 400
rect 53088 0 53144 400
rect 53368 0 53424 400
rect 53648 0 53704 400
rect 53928 0 53984 400
rect 54208 0 54264 400
rect 54488 0 54544 400
rect 54768 0 54824 400
rect 55048 0 55104 400
rect 55328 0 55384 400
rect 55608 0 55664 400
rect 55888 0 55944 400
rect 56168 0 56224 400
rect 56448 0 56504 400
rect 56728 0 56784 400
rect 57008 0 57064 400
rect 57288 0 57344 400
rect 57568 0 57624 400
rect 57848 0 57904 400
rect 58128 0 58184 400
rect 58408 0 58464 400
rect 58688 0 58744 400
rect 58968 0 59024 400
rect 59248 0 59304 400
rect 59528 0 59584 400
rect 59808 0 59864 400
rect 60088 0 60144 400
rect 60368 0 60424 400
rect 60648 0 60704 400
rect 60928 0 60984 400
rect 61208 0 61264 400
rect 61488 0 61544 400
rect 61768 0 61824 400
rect 62048 0 62104 400
rect 62328 0 62384 400
rect 62608 0 62664 400
rect 62888 0 62944 400
rect 63168 0 63224 400
rect 63448 0 63504 400
rect 63728 0 63784 400
rect 64008 0 64064 400
rect 64288 0 64344 400
rect 64568 0 64624 400
rect 64848 0 64904 400
rect 65128 0 65184 400
rect 65408 0 65464 400
rect 65688 0 65744 400
rect 65968 0 66024 400
rect 66248 0 66304 400
rect 66528 0 66584 400
rect 66808 0 66864 400
rect 67088 0 67144 400
rect 67368 0 67424 400
rect 67648 0 67704 400
rect 67928 0 67984 400
rect 68208 0 68264 400
rect 68488 0 68544 400
rect 68768 0 68824 400
rect 69048 0 69104 400
rect 69328 0 69384 400
rect 69608 0 69664 400
rect 69888 0 69944 400
rect 70168 0 70224 400
rect 70448 0 70504 400
rect 70728 0 70784 400
rect 71008 0 71064 400
rect 71288 0 71344 400
rect 71568 0 71624 400
rect 71848 0 71904 400
rect 72128 0 72184 400
rect 72408 0 72464 400
rect 72688 0 72744 400
rect 72968 0 73024 400
rect 73248 0 73304 400
rect 73528 0 73584 400
rect 73808 0 73864 400
rect 74088 0 74144 400
rect 74368 0 74424 400
rect 74648 0 74704 400
rect 74928 0 74984 400
rect 75208 0 75264 400
rect 75488 0 75544 400
rect 75768 0 75824 400
rect 76048 0 76104 400
rect 76328 0 76384 400
rect 76608 0 76664 400
rect 76888 0 76944 400
rect 77168 0 77224 400
rect 77448 0 77504 400
rect 77728 0 77784 400
rect 78008 0 78064 400
rect 78288 0 78344 400
rect 78568 0 78624 400
rect 78848 0 78904 400
rect 79128 0 79184 400
rect 79408 0 79464 400
rect 79688 0 79744 400
rect 79968 0 80024 400
rect 80248 0 80304 400
rect 80528 0 80584 400
rect 80808 0 80864 400
rect 81088 0 81144 400
rect 81368 0 81424 400
rect 81648 0 81704 400
rect 81928 0 81984 400
rect 82208 0 82264 400
rect 82488 0 82544 400
rect 82768 0 82824 400
rect 83048 0 83104 400
rect 83328 0 83384 400
rect 83608 0 83664 400
rect 83888 0 83944 400
rect 84168 0 84224 400
rect 84448 0 84504 400
rect 84728 0 84784 400
rect 85008 0 85064 400
rect 85288 0 85344 400
rect 85568 0 85624 400
rect 85848 0 85904 400
rect 86128 0 86184 400
rect 86408 0 86464 400
rect 86688 0 86744 400
rect 86968 0 87024 400
rect 87248 0 87304 400
rect 87528 0 87584 400
rect 87808 0 87864 400
rect 88088 0 88144 400
rect 88368 0 88424 400
rect 88648 0 88704 400
rect 88928 0 88984 400
rect 89208 0 89264 400
rect 89488 0 89544 400
rect 89768 0 89824 400
rect 90048 0 90104 400
rect 90328 0 90384 400
rect 90608 0 90664 400
rect 90888 0 90944 400
rect 91168 0 91224 400
rect 91448 0 91504 400
rect 91728 0 91784 400
rect 92008 0 92064 400
rect 92288 0 92344 400
rect 92568 0 92624 400
rect 92848 0 92904 400
rect 93128 0 93184 400
rect 93408 0 93464 400
rect 93688 0 93744 400
rect 93968 0 94024 400
rect 94248 0 94304 400
rect 94528 0 94584 400
rect 94808 0 94864 400
rect 95088 0 95144 400
rect 95368 0 95424 400
rect 95648 0 95704 400
rect 95928 0 95984 400
rect 96208 0 96264 400
rect 96488 0 96544 400
rect 96768 0 96824 400
rect 97048 0 97104 400
rect 97328 0 97384 400
rect 97608 0 97664 400
rect 97888 0 97944 400
rect 98168 0 98224 400
rect 98448 0 98504 400
rect 98728 0 98784 400
rect 99008 0 99064 400
rect 99288 0 99344 400
rect 99568 0 99624 400
rect 99848 0 99904 400
rect 100128 0 100184 400
rect 100408 0 100464 400
rect 100688 0 100744 400
rect 100968 0 101024 400
rect 101248 0 101304 400
rect 101528 0 101584 400
rect 101808 0 101864 400
rect 102088 0 102144 400
rect 102368 0 102424 400
rect 102648 0 102704 400
rect 102928 0 102984 400
rect 103208 0 103264 400
rect 103488 0 103544 400
rect 103768 0 103824 400
rect 104048 0 104104 400
rect 104328 0 104384 400
rect 104608 0 104664 400
rect 104888 0 104944 400
rect 105168 0 105224 400
rect 105448 0 105504 400
rect 105728 0 105784 400
rect 106008 0 106064 400
rect 106288 0 106344 400
rect 106568 0 106624 400
rect 106848 0 106904 400
rect 107128 0 107184 400
rect 107408 0 107464 400
rect 107688 0 107744 400
rect 107968 0 108024 400
rect 108248 0 108304 400
rect 108528 0 108584 400
rect 108808 0 108864 400
rect 109088 0 109144 400
rect 109368 0 109424 400
rect 109648 0 109704 400
rect 109928 0 109984 400
rect 110208 0 110264 400
rect 110488 0 110544 400
rect 110768 0 110824 400
rect 111048 0 111104 400
rect 111328 0 111384 400
rect 111608 0 111664 400
rect 111888 0 111944 400
rect 112168 0 112224 400
rect 112448 0 112504 400
rect 112728 0 112784 400
rect 113008 0 113064 400
rect 113288 0 113344 400
rect 113568 0 113624 400
rect 113848 0 113904 400
rect 114128 0 114184 400
rect 114408 0 114464 400
rect 114688 0 114744 400
rect 114968 0 115024 400
rect 115248 0 115304 400
rect 115528 0 115584 400
rect 115808 0 115864 400
rect 116088 0 116144 400
rect 116368 0 116424 400
rect 116648 0 116704 400
rect 116928 0 116984 400
rect 117208 0 117264 400
rect 117488 0 117544 400
rect 117768 0 117824 400
rect 118048 0 118104 400
rect 118328 0 118384 400
rect 118608 0 118664 400
rect 118888 0 118944 400
rect 119168 0 119224 400
rect 119448 0 119504 400
rect 119728 0 119784 400
rect 120008 0 120064 400
rect 120288 0 120344 400
rect 120568 0 120624 400
rect 120848 0 120904 400
rect 121128 0 121184 400
rect 121408 0 121464 400
rect 121688 0 121744 400
rect 121968 0 122024 400
rect 122248 0 122304 400
rect 122528 0 122584 400
rect 122808 0 122864 400
rect 123088 0 123144 400
rect 123368 0 123424 400
rect 123648 0 123704 400
rect 123928 0 123984 400
rect 124208 0 124264 400
rect 124488 0 124544 400
rect 124768 0 124824 400
rect 125048 0 125104 400
rect 125328 0 125384 400
rect 125608 0 125664 400
rect 125888 0 125944 400
rect 126168 0 126224 400
rect 126448 0 126504 400
rect 126728 0 126784 400
rect 127008 0 127064 400
rect 127288 0 127344 400
rect 127568 0 127624 400
rect 127848 0 127904 400
rect 128128 0 128184 400
rect 128408 0 128464 400
rect 128688 0 128744 400
rect 128968 0 129024 400
rect 129248 0 129304 400
rect 129528 0 129584 400
rect 129808 0 129864 400
rect 130088 0 130144 400
rect 130368 0 130424 400
rect 130648 0 130704 400
rect 130928 0 130984 400
rect 131208 0 131264 400
rect 131488 0 131544 400
rect 131768 0 131824 400
rect 132048 0 132104 400
rect 132328 0 132384 400
rect 132608 0 132664 400
rect 132888 0 132944 400
rect 133168 0 133224 400
rect 133448 0 133504 400
rect 133728 0 133784 400
rect 134008 0 134064 400
rect 134288 0 134344 400
rect 134568 0 134624 400
rect 134848 0 134904 400
rect 135128 0 135184 400
rect 135408 0 135464 400
rect 135688 0 135744 400
rect 135968 0 136024 400
rect 136248 0 136304 400
rect 136528 0 136584 400
rect 136808 0 136864 400
rect 137088 0 137144 400
rect 137368 0 137424 400
rect 137648 0 137704 400
rect 137928 0 137984 400
rect 138208 0 138264 400
rect 138488 0 138544 400
rect 138768 0 138824 400
rect 139048 0 139104 400
rect 139328 0 139384 400
rect 139608 0 139664 400
rect 139888 0 139944 400
rect 140168 0 140224 400
rect 140448 0 140504 400
rect 140728 0 140784 400
rect 141008 0 141064 400
rect 141288 0 141344 400
rect 141568 0 141624 400
rect 141848 0 141904 400
rect 142128 0 142184 400
rect 142408 0 142464 400
rect 142688 0 142744 400
rect 142968 0 143024 400
rect 143248 0 143304 400
rect 143528 0 143584 400
rect 143808 0 143864 400
<< obsm2 >>
rect 910 149570 2154 149600
rect 2270 149570 3442 149600
rect 3558 149570 4730 149600
rect 4846 149570 6018 149600
rect 6134 149570 7306 149600
rect 7422 149570 8594 149600
rect 8710 149570 9882 149600
rect 9998 149570 11170 149600
rect 11286 149570 12458 149600
rect 12574 149570 13746 149600
rect 13862 149570 15034 149600
rect 15150 149570 16322 149600
rect 16438 149570 17610 149600
rect 17726 149570 18898 149600
rect 19014 149570 20186 149600
rect 20302 149570 21474 149600
rect 21590 149570 22762 149600
rect 22878 149570 24050 149600
rect 24166 149570 25338 149600
rect 25454 149570 26626 149600
rect 26742 149570 27914 149600
rect 28030 149570 29202 149600
rect 29318 149570 30490 149600
rect 30606 149570 31778 149600
rect 31894 149570 33066 149600
rect 33182 149570 34354 149600
rect 34470 149570 35642 149600
rect 35758 149570 36930 149600
rect 37046 149570 38218 149600
rect 38334 149570 39506 149600
rect 39622 149570 40794 149600
rect 40910 149570 42082 149600
rect 42198 149570 43370 149600
rect 43486 149570 44658 149600
rect 44774 149570 45946 149600
rect 46062 149570 47234 149600
rect 47350 149570 48522 149600
rect 48638 149570 49810 149600
rect 49926 149570 51098 149600
rect 51214 149570 52386 149600
rect 52502 149570 53674 149600
rect 53790 149570 54962 149600
rect 55078 149570 56250 149600
rect 56366 149570 57538 149600
rect 57654 149570 58826 149600
rect 58942 149570 60114 149600
rect 60230 149570 61402 149600
rect 61518 149570 62690 149600
rect 62806 149570 63978 149600
rect 64094 149570 65266 149600
rect 65382 149570 66554 149600
rect 66670 149570 67842 149600
rect 67958 149570 69130 149600
rect 69246 149570 70418 149600
rect 70534 149570 71706 149600
rect 71822 149570 72994 149600
rect 73110 149570 74282 149600
rect 74398 149570 75570 149600
rect 75686 149570 76858 149600
rect 76974 149570 78146 149600
rect 78262 149570 79434 149600
rect 79550 149570 80722 149600
rect 80838 149570 82010 149600
rect 82126 149570 83298 149600
rect 83414 149570 84586 149600
rect 84702 149570 85874 149600
rect 85990 149570 87162 149600
rect 87278 149570 88450 149600
rect 88566 149570 89738 149600
rect 89854 149570 91026 149600
rect 91142 149570 92314 149600
rect 92430 149570 93602 149600
rect 93718 149570 94890 149600
rect 95006 149570 96178 149600
rect 96294 149570 97466 149600
rect 97582 149570 98754 149600
rect 98870 149570 100042 149600
rect 100158 149570 101330 149600
rect 101446 149570 102618 149600
rect 102734 149570 103906 149600
rect 104022 149570 105194 149600
rect 105310 149570 106482 149600
rect 106598 149570 107770 149600
rect 107886 149570 109058 149600
rect 109174 149570 110346 149600
rect 110462 149570 111634 149600
rect 111750 149570 112922 149600
rect 113038 149570 114210 149600
rect 114326 149570 115498 149600
rect 115614 149570 116786 149600
rect 116902 149570 118074 149600
rect 118190 149570 119362 149600
rect 119478 149570 120650 149600
rect 120766 149570 121938 149600
rect 122054 149570 123226 149600
rect 123342 149570 124514 149600
rect 124630 149570 125802 149600
rect 125918 149570 127090 149600
rect 127206 149570 128378 149600
rect 128494 149570 129666 149600
rect 129782 149570 130954 149600
rect 131070 149570 132242 149600
rect 132358 149570 133530 149600
rect 133646 149570 134818 149600
rect 134934 149570 136106 149600
rect 136222 149570 137394 149600
rect 137510 149570 138682 149600
rect 138798 149570 139970 149600
rect 140086 149570 141258 149600
rect 141374 149570 142546 149600
rect 142662 149570 143834 149600
rect 143950 149570 145122 149600
rect 145238 149570 146410 149600
rect 146526 149570 147698 149600
rect 147814 149570 149058 149600
rect 910 430 149058 149570
rect 910 400 6018 430
rect 6134 400 6298 430
rect 6414 400 6578 430
rect 6694 400 6858 430
rect 6974 400 7138 430
rect 7254 400 7418 430
rect 7534 400 7698 430
rect 7814 400 7978 430
rect 8094 400 8258 430
rect 8374 400 8538 430
rect 8654 400 8818 430
rect 8934 400 9098 430
rect 9214 400 9378 430
rect 9494 400 9658 430
rect 9774 400 9938 430
rect 10054 400 10218 430
rect 10334 400 10498 430
rect 10614 400 10778 430
rect 10894 400 11058 430
rect 11174 400 11338 430
rect 11454 400 11618 430
rect 11734 400 11898 430
rect 12014 400 12178 430
rect 12294 400 12458 430
rect 12574 400 12738 430
rect 12854 400 13018 430
rect 13134 400 13298 430
rect 13414 400 13578 430
rect 13694 400 13858 430
rect 13974 400 14138 430
rect 14254 400 14418 430
rect 14534 400 14698 430
rect 14814 400 14978 430
rect 15094 400 15258 430
rect 15374 400 15538 430
rect 15654 400 15818 430
rect 15934 400 16098 430
rect 16214 400 16378 430
rect 16494 400 16658 430
rect 16774 400 16938 430
rect 17054 400 17218 430
rect 17334 400 17498 430
rect 17614 400 17778 430
rect 17894 400 18058 430
rect 18174 400 18338 430
rect 18454 400 18618 430
rect 18734 400 18898 430
rect 19014 400 19178 430
rect 19294 400 19458 430
rect 19574 400 19738 430
rect 19854 400 20018 430
rect 20134 400 20298 430
rect 20414 400 20578 430
rect 20694 400 20858 430
rect 20974 400 21138 430
rect 21254 400 21418 430
rect 21534 400 21698 430
rect 21814 400 21978 430
rect 22094 400 22258 430
rect 22374 400 22538 430
rect 22654 400 22818 430
rect 22934 400 23098 430
rect 23214 400 23378 430
rect 23494 400 23658 430
rect 23774 400 23938 430
rect 24054 400 24218 430
rect 24334 400 24498 430
rect 24614 400 24778 430
rect 24894 400 25058 430
rect 25174 400 25338 430
rect 25454 400 25618 430
rect 25734 400 25898 430
rect 26014 400 26178 430
rect 26294 400 26458 430
rect 26574 400 26738 430
rect 26854 400 27018 430
rect 27134 400 27298 430
rect 27414 400 27578 430
rect 27694 400 27858 430
rect 27974 400 28138 430
rect 28254 400 28418 430
rect 28534 400 28698 430
rect 28814 400 28978 430
rect 29094 400 29258 430
rect 29374 400 29538 430
rect 29654 400 29818 430
rect 29934 400 30098 430
rect 30214 400 30378 430
rect 30494 400 30658 430
rect 30774 400 30938 430
rect 31054 400 31218 430
rect 31334 400 31498 430
rect 31614 400 31778 430
rect 31894 400 32058 430
rect 32174 400 32338 430
rect 32454 400 32618 430
rect 32734 400 32898 430
rect 33014 400 33178 430
rect 33294 400 33458 430
rect 33574 400 33738 430
rect 33854 400 34018 430
rect 34134 400 34298 430
rect 34414 400 34578 430
rect 34694 400 34858 430
rect 34974 400 35138 430
rect 35254 400 35418 430
rect 35534 400 35698 430
rect 35814 400 35978 430
rect 36094 400 36258 430
rect 36374 400 36538 430
rect 36654 400 36818 430
rect 36934 400 37098 430
rect 37214 400 37378 430
rect 37494 400 37658 430
rect 37774 400 37938 430
rect 38054 400 38218 430
rect 38334 400 38498 430
rect 38614 400 38778 430
rect 38894 400 39058 430
rect 39174 400 39338 430
rect 39454 400 39618 430
rect 39734 400 39898 430
rect 40014 400 40178 430
rect 40294 400 40458 430
rect 40574 400 40738 430
rect 40854 400 41018 430
rect 41134 400 41298 430
rect 41414 400 41578 430
rect 41694 400 41858 430
rect 41974 400 42138 430
rect 42254 400 42418 430
rect 42534 400 42698 430
rect 42814 400 42978 430
rect 43094 400 43258 430
rect 43374 400 43538 430
rect 43654 400 43818 430
rect 43934 400 44098 430
rect 44214 400 44378 430
rect 44494 400 44658 430
rect 44774 400 44938 430
rect 45054 400 45218 430
rect 45334 400 45498 430
rect 45614 400 45778 430
rect 45894 400 46058 430
rect 46174 400 46338 430
rect 46454 400 46618 430
rect 46734 400 46898 430
rect 47014 400 47178 430
rect 47294 400 47458 430
rect 47574 400 47738 430
rect 47854 400 48018 430
rect 48134 400 48298 430
rect 48414 400 48578 430
rect 48694 400 48858 430
rect 48974 400 49138 430
rect 49254 400 49418 430
rect 49534 400 49698 430
rect 49814 400 49978 430
rect 50094 400 50258 430
rect 50374 400 50538 430
rect 50654 400 50818 430
rect 50934 400 51098 430
rect 51214 400 51378 430
rect 51494 400 51658 430
rect 51774 400 51938 430
rect 52054 400 52218 430
rect 52334 400 52498 430
rect 52614 400 52778 430
rect 52894 400 53058 430
rect 53174 400 53338 430
rect 53454 400 53618 430
rect 53734 400 53898 430
rect 54014 400 54178 430
rect 54294 400 54458 430
rect 54574 400 54738 430
rect 54854 400 55018 430
rect 55134 400 55298 430
rect 55414 400 55578 430
rect 55694 400 55858 430
rect 55974 400 56138 430
rect 56254 400 56418 430
rect 56534 400 56698 430
rect 56814 400 56978 430
rect 57094 400 57258 430
rect 57374 400 57538 430
rect 57654 400 57818 430
rect 57934 400 58098 430
rect 58214 400 58378 430
rect 58494 400 58658 430
rect 58774 400 58938 430
rect 59054 400 59218 430
rect 59334 400 59498 430
rect 59614 400 59778 430
rect 59894 400 60058 430
rect 60174 400 60338 430
rect 60454 400 60618 430
rect 60734 400 60898 430
rect 61014 400 61178 430
rect 61294 400 61458 430
rect 61574 400 61738 430
rect 61854 400 62018 430
rect 62134 400 62298 430
rect 62414 400 62578 430
rect 62694 400 62858 430
rect 62974 400 63138 430
rect 63254 400 63418 430
rect 63534 400 63698 430
rect 63814 400 63978 430
rect 64094 400 64258 430
rect 64374 400 64538 430
rect 64654 400 64818 430
rect 64934 400 65098 430
rect 65214 400 65378 430
rect 65494 400 65658 430
rect 65774 400 65938 430
rect 66054 400 66218 430
rect 66334 400 66498 430
rect 66614 400 66778 430
rect 66894 400 67058 430
rect 67174 400 67338 430
rect 67454 400 67618 430
rect 67734 400 67898 430
rect 68014 400 68178 430
rect 68294 400 68458 430
rect 68574 400 68738 430
rect 68854 400 69018 430
rect 69134 400 69298 430
rect 69414 400 69578 430
rect 69694 400 69858 430
rect 69974 400 70138 430
rect 70254 400 70418 430
rect 70534 400 70698 430
rect 70814 400 70978 430
rect 71094 400 71258 430
rect 71374 400 71538 430
rect 71654 400 71818 430
rect 71934 400 72098 430
rect 72214 400 72378 430
rect 72494 400 72658 430
rect 72774 400 72938 430
rect 73054 400 73218 430
rect 73334 400 73498 430
rect 73614 400 73778 430
rect 73894 400 74058 430
rect 74174 400 74338 430
rect 74454 400 74618 430
rect 74734 400 74898 430
rect 75014 400 75178 430
rect 75294 400 75458 430
rect 75574 400 75738 430
rect 75854 400 76018 430
rect 76134 400 76298 430
rect 76414 400 76578 430
rect 76694 400 76858 430
rect 76974 400 77138 430
rect 77254 400 77418 430
rect 77534 400 77698 430
rect 77814 400 77978 430
rect 78094 400 78258 430
rect 78374 400 78538 430
rect 78654 400 78818 430
rect 78934 400 79098 430
rect 79214 400 79378 430
rect 79494 400 79658 430
rect 79774 400 79938 430
rect 80054 400 80218 430
rect 80334 400 80498 430
rect 80614 400 80778 430
rect 80894 400 81058 430
rect 81174 400 81338 430
rect 81454 400 81618 430
rect 81734 400 81898 430
rect 82014 400 82178 430
rect 82294 400 82458 430
rect 82574 400 82738 430
rect 82854 400 83018 430
rect 83134 400 83298 430
rect 83414 400 83578 430
rect 83694 400 83858 430
rect 83974 400 84138 430
rect 84254 400 84418 430
rect 84534 400 84698 430
rect 84814 400 84978 430
rect 85094 400 85258 430
rect 85374 400 85538 430
rect 85654 400 85818 430
rect 85934 400 86098 430
rect 86214 400 86378 430
rect 86494 400 86658 430
rect 86774 400 86938 430
rect 87054 400 87218 430
rect 87334 400 87498 430
rect 87614 400 87778 430
rect 87894 400 88058 430
rect 88174 400 88338 430
rect 88454 400 88618 430
rect 88734 400 88898 430
rect 89014 400 89178 430
rect 89294 400 89458 430
rect 89574 400 89738 430
rect 89854 400 90018 430
rect 90134 400 90298 430
rect 90414 400 90578 430
rect 90694 400 90858 430
rect 90974 400 91138 430
rect 91254 400 91418 430
rect 91534 400 91698 430
rect 91814 400 91978 430
rect 92094 400 92258 430
rect 92374 400 92538 430
rect 92654 400 92818 430
rect 92934 400 93098 430
rect 93214 400 93378 430
rect 93494 400 93658 430
rect 93774 400 93938 430
rect 94054 400 94218 430
rect 94334 400 94498 430
rect 94614 400 94778 430
rect 94894 400 95058 430
rect 95174 400 95338 430
rect 95454 400 95618 430
rect 95734 400 95898 430
rect 96014 400 96178 430
rect 96294 400 96458 430
rect 96574 400 96738 430
rect 96854 400 97018 430
rect 97134 400 97298 430
rect 97414 400 97578 430
rect 97694 400 97858 430
rect 97974 400 98138 430
rect 98254 400 98418 430
rect 98534 400 98698 430
rect 98814 400 98978 430
rect 99094 400 99258 430
rect 99374 400 99538 430
rect 99654 400 99818 430
rect 99934 400 100098 430
rect 100214 400 100378 430
rect 100494 400 100658 430
rect 100774 400 100938 430
rect 101054 400 101218 430
rect 101334 400 101498 430
rect 101614 400 101778 430
rect 101894 400 102058 430
rect 102174 400 102338 430
rect 102454 400 102618 430
rect 102734 400 102898 430
rect 103014 400 103178 430
rect 103294 400 103458 430
rect 103574 400 103738 430
rect 103854 400 104018 430
rect 104134 400 104298 430
rect 104414 400 104578 430
rect 104694 400 104858 430
rect 104974 400 105138 430
rect 105254 400 105418 430
rect 105534 400 105698 430
rect 105814 400 105978 430
rect 106094 400 106258 430
rect 106374 400 106538 430
rect 106654 400 106818 430
rect 106934 400 107098 430
rect 107214 400 107378 430
rect 107494 400 107658 430
rect 107774 400 107938 430
rect 108054 400 108218 430
rect 108334 400 108498 430
rect 108614 400 108778 430
rect 108894 400 109058 430
rect 109174 400 109338 430
rect 109454 400 109618 430
rect 109734 400 109898 430
rect 110014 400 110178 430
rect 110294 400 110458 430
rect 110574 400 110738 430
rect 110854 400 111018 430
rect 111134 400 111298 430
rect 111414 400 111578 430
rect 111694 400 111858 430
rect 111974 400 112138 430
rect 112254 400 112418 430
rect 112534 400 112698 430
rect 112814 400 112978 430
rect 113094 400 113258 430
rect 113374 400 113538 430
rect 113654 400 113818 430
rect 113934 400 114098 430
rect 114214 400 114378 430
rect 114494 400 114658 430
rect 114774 400 114938 430
rect 115054 400 115218 430
rect 115334 400 115498 430
rect 115614 400 115778 430
rect 115894 400 116058 430
rect 116174 400 116338 430
rect 116454 400 116618 430
rect 116734 400 116898 430
rect 117014 400 117178 430
rect 117294 400 117458 430
rect 117574 400 117738 430
rect 117854 400 118018 430
rect 118134 400 118298 430
rect 118414 400 118578 430
rect 118694 400 118858 430
rect 118974 400 119138 430
rect 119254 400 119418 430
rect 119534 400 119698 430
rect 119814 400 119978 430
rect 120094 400 120258 430
rect 120374 400 120538 430
rect 120654 400 120818 430
rect 120934 400 121098 430
rect 121214 400 121378 430
rect 121494 400 121658 430
rect 121774 400 121938 430
rect 122054 400 122218 430
rect 122334 400 122498 430
rect 122614 400 122778 430
rect 122894 400 123058 430
rect 123174 400 123338 430
rect 123454 400 123618 430
rect 123734 400 123898 430
rect 124014 400 124178 430
rect 124294 400 124458 430
rect 124574 400 124738 430
rect 124854 400 125018 430
rect 125134 400 125298 430
rect 125414 400 125578 430
rect 125694 400 125858 430
rect 125974 400 126138 430
rect 126254 400 126418 430
rect 126534 400 126698 430
rect 126814 400 126978 430
rect 127094 400 127258 430
rect 127374 400 127538 430
rect 127654 400 127818 430
rect 127934 400 128098 430
rect 128214 400 128378 430
rect 128494 400 128658 430
rect 128774 400 128938 430
rect 129054 400 129218 430
rect 129334 400 129498 430
rect 129614 400 129778 430
rect 129894 400 130058 430
rect 130174 400 130338 430
rect 130454 400 130618 430
rect 130734 400 130898 430
rect 131014 400 131178 430
rect 131294 400 131458 430
rect 131574 400 131738 430
rect 131854 400 132018 430
rect 132134 400 132298 430
rect 132414 400 132578 430
rect 132694 400 132858 430
rect 132974 400 133138 430
rect 133254 400 133418 430
rect 133534 400 133698 430
rect 133814 400 133978 430
rect 134094 400 134258 430
rect 134374 400 134538 430
rect 134654 400 134818 430
rect 134934 400 135098 430
rect 135214 400 135378 430
rect 135494 400 135658 430
rect 135774 400 135938 430
rect 136054 400 136218 430
rect 136334 400 136498 430
rect 136614 400 136778 430
rect 136894 400 137058 430
rect 137174 400 137338 430
rect 137454 400 137618 430
rect 137734 400 137898 430
rect 138014 400 138178 430
rect 138294 400 138458 430
rect 138574 400 138738 430
rect 138854 400 139018 430
rect 139134 400 139298 430
rect 139414 400 139578 430
rect 139694 400 139858 430
rect 139974 400 140138 430
rect 140254 400 140418 430
rect 140534 400 140698 430
rect 140814 400 140978 430
rect 141094 400 141258 430
rect 141374 400 141538 430
rect 141654 400 141818 430
rect 141934 400 142098 430
rect 142214 400 142378 430
rect 142494 400 142658 430
rect 142774 400 142938 430
rect 143054 400 143218 430
rect 143334 400 143498 430
rect 143614 400 143778 430
rect 143894 400 149058 430
<< obsm3 >>
rect 905 1554 149063 148190
<< metal4 >>
rect 2224 1538 2384 148206
rect 9904 1538 10064 148206
rect 17584 1538 17744 148206
rect 25264 1538 25424 148206
rect 32944 1538 33104 148206
rect 40624 1538 40784 148206
rect 48304 1538 48464 148206
rect 55984 1538 56144 148206
rect 63664 1538 63824 148206
rect 71344 1538 71504 148206
rect 79024 1538 79184 148206
rect 86704 1538 86864 148206
rect 94384 1538 94544 148206
rect 102064 1538 102224 148206
rect 109744 1538 109904 148206
rect 117424 1538 117584 148206
rect 125104 1538 125264 148206
rect 132784 1538 132944 148206
rect 140464 1538 140624 148206
rect 148144 1538 148304 148206
<< obsm4 >>
rect 2142 2641 2194 147999
rect 2414 2641 9874 147999
rect 10094 2641 17554 147999
rect 17774 2641 25234 147999
rect 25454 2641 32914 147999
rect 33134 2641 40594 147999
rect 40814 2641 48274 147999
rect 48494 2641 55954 147999
rect 56174 2641 63634 147999
rect 63854 2641 71314 147999
rect 71534 2641 78994 147999
rect 79214 2641 86674 147999
rect 86894 2641 94354 147999
rect 94574 2641 102034 147999
rect 102254 2641 109714 147999
rect 109934 2641 117394 147999
rect 117614 2641 125074 147999
rect 125294 2641 132754 147999
rect 132974 2641 140434 147999
rect 140654 2641 148050 147999
<< obsm5 >>
rect 2134 3758 147050 140722
<< labels >>
rlabel metal2 s 2184 149600 2240 150000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 40824 149600 40880 150000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 44688 149600 44744 150000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 48552 149600 48608 150000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 52416 149600 52472 150000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 56280 149600 56336 150000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 60144 149600 60200 150000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 64008 149600 64064 150000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 67872 149600 67928 150000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 71736 149600 71792 150000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 75600 149600 75656 150000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6048 149600 6104 150000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 79464 149600 79520 150000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 83328 149600 83384 150000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 87192 149600 87248 150000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 91056 149600 91112 150000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 94920 149600 94976 150000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 98784 149600 98840 150000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 102648 149600 102704 150000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 106512 149600 106568 150000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 110376 149600 110432 150000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 114240 149600 114296 150000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9912 149600 9968 150000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 118104 149600 118160 150000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 121968 149600 122024 150000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 125832 149600 125888 150000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 129696 149600 129752 150000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 133560 149600 133616 150000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 137424 149600 137480 150000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 141288 149600 141344 150000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 145152 149600 145208 150000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13776 149600 13832 150000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17640 149600 17696 150000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21504 149600 21560 150000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 25368 149600 25424 150000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 29232 149600 29288 150000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 33096 149600 33152 150000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 36960 149600 37016 150000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3472 149600 3528 150000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 42112 149600 42168 150000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 45976 149600 46032 150000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 49840 149600 49896 150000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 53704 149600 53760 150000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 57568 149600 57624 150000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 61432 149600 61488 150000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 65296 149600 65352 150000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 69160 149600 69216 150000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 73024 149600 73080 150000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 76888 149600 76944 150000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7336 149600 7392 150000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 80752 149600 80808 150000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 84616 149600 84672 150000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 88480 149600 88536 150000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 92344 149600 92400 150000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 96208 149600 96264 150000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 100072 149600 100128 150000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 103936 149600 103992 150000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 107800 149600 107856 150000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 111664 149600 111720 150000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 115528 149600 115584 150000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11200 149600 11256 150000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 119392 149600 119448 150000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 123256 149600 123312 150000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 127120 149600 127176 150000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 130984 149600 131040 150000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 134848 149600 134904 150000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 138712 149600 138768 150000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 142576 149600 142632 150000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 146440 149600 146496 150000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15064 149600 15120 150000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 18928 149600 18984 150000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 22792 149600 22848 150000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 26656 149600 26712 150000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 30520 149600 30576 150000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 34384 149600 34440 150000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 38248 149600 38304 150000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4760 149600 4816 150000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 43400 149600 43456 150000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 47264 149600 47320 150000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 51128 149600 51184 150000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 54992 149600 55048 150000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 58856 149600 58912 150000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 62720 149600 62776 150000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 66584 149600 66640 150000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 70448 149600 70504 150000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 74312 149600 74368 150000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 78176 149600 78232 150000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8624 149600 8680 150000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 82040 149600 82096 150000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 85904 149600 85960 150000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 89768 149600 89824 150000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 93632 149600 93688 150000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 97496 149600 97552 150000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 101360 149600 101416 150000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 105224 149600 105280 150000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 109088 149600 109144 150000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 112952 149600 113008 150000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 116816 149600 116872 150000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12488 149600 12544 150000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 120680 149600 120736 150000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 124544 149600 124600 150000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 128408 149600 128464 150000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 132272 149600 132328 150000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 136136 149600 136192 150000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 140000 149600 140056 150000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 143864 149600 143920 150000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 147728 149600 147784 150000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16352 149600 16408 150000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20216 149600 20272 150000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24080 149600 24136 150000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 27944 149600 28000 150000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 31808 149600 31864 150000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 35672 149600 35728 150000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 39536 149600 39592 150000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 143248 0 143304 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 143528 0 143584 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 143808 0 143864 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 119728 0 119784 400 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 120568 0 120624 400 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 121408 0 121464 400 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 122248 0 122304 400 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 123088 0 123144 400 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 123928 0 123984 400 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 124768 0 124824 400 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 125608 0 125664 400 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 127288 0 127344 400 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 128128 0 128184 400 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 128968 0 129024 400 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 129808 0 129864 400 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 130648 0 130704 400 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 131488 0 131544 400 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 132328 0 132384 400 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 133168 0 133224 400 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 134008 0 134064 400 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 134848 0 134904 400 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 135688 0 135744 400 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 136528 0 136584 400 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 137368 0 137424 400 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 138208 0 138264 400 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 139048 0 139104 400 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 140728 0 140784 400 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 141568 0 141624 400 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 142408 0 142464 400 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 46648 0 46704 400 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 48328 0 48384 400 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 51688 0 51744 400 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 36568 0 36624 400 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 53368 0 53424 400 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 55048 0 55104 400 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 56728 0 56784 400 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 58408 0 58464 400 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 60088 0 60144 400 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 61768 0 61824 400 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 62608 0 62664 400 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 63448 0 63504 400 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 65128 0 65184 400 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 66808 0 66864 400 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 68488 0 68544 400 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 38248 0 38304 400 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 70168 0 70224 400 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 71848 0 71904 400 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 73528 0 73584 400 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 75208 0 75264 400 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 76048 0 76104 400 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 76888 0 76944 400 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 78568 0 78624 400 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 80248 0 80304 400 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 81928 0 81984 400 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 82768 0 82824 400 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 83608 0 83664 400 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 86968 0 87024 400 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 87808 0 87864 400 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 88648 0 88704 400 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 89488 0 89544 400 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 90328 0 90384 400 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 91168 0 91224 400 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 92008 0 92064 400 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 93688 0 93744 400 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 94528 0 94584 400 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 95368 0 95424 400 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 97048 0 97104 400 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 97888 0 97944 400 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 98728 0 98784 400 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 99568 0 99624 400 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 100408 0 100464 400 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 101248 0 101304 400 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 102088 0 102144 400 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 41608 0 41664 400 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 102928 0 102984 400 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 103768 0 103824 400 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 104608 0 104664 400 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 105448 0 105504 400 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 106288 0 106344 400 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 107128 0 107184 400 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 107968 0 108024 400 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 108808 0 108864 400 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 109648 0 109704 400 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 110488 0 110544 400 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 111328 0 111384 400 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 112168 0 112224 400 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 113848 0 113904 400 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 114688 0 114744 400 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 115528 0 115584 400 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 116368 0 116424 400 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 117208 0 117264 400 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 118048 0 118104 400 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 118888 0 118944 400 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43288 0 43344 400 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 36008 0 36064 400 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 120008 0 120064 400 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 120848 0 120904 400 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 121688 0 121744 400 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 122528 0 122584 400 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 123368 0 123424 400 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 124208 0 124264 400 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 125048 0 125104 400 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 125888 0 125944 400 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 126728 0 126784 400 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 127568 0 127624 400 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 44408 0 44464 400 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 128408 0 128464 400 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 129248 0 129304 400 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 130088 0 130144 400 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 131768 0 131824 400 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 132608 0 132664 400 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 133448 0 133504 400 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 134288 0 134344 400 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 135128 0 135184 400 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 135968 0 136024 400 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 45248 0 45304 400 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 136808 0 136864 400 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 137648 0 137704 400 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 138488 0 138544 400 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 139328 0 139384 400 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 140168 0 140224 400 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 141008 0 141064 400 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 141848 0 141904 400 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 142688 0 142744 400 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 46088 0 46144 400 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 46928 0 46984 400 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 47768 0 47824 400 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 48608 0 48664 400 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 49448 0 49504 400 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 50288 0 50344 400 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 51128 0 51184 400 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 36848 0 36904 400 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 52808 0 52864 400 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 53648 0 53704 400 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 54488 0 54544 400 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 55328 0 55384 400 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 56168 0 56224 400 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 57848 0 57904 400 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 58688 0 58744 400 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 59528 0 59584 400 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 60368 0 60424 400 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 37688 0 37744 400 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 61208 0 61264 400 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 62048 0 62104 400 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 62888 0 62944 400 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 64568 0 64624 400 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 65408 0 65464 400 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 66248 0 66304 400 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 67088 0 67144 400 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 67928 0 67984 400 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 38528 0 38584 400 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 69608 0 69664 400 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 70448 0 70504 400 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 71288 0 71344 400 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 72128 0 72184 400 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 72968 0 73024 400 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 73808 0 73864 400 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 74648 0 74704 400 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 75488 0 75544 400 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 76328 0 76384 400 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 39368 0 39424 400 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 78008 0 78064 400 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 78848 0 78904 400 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 79688 0 79744 400 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 80528 0 80584 400 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 81368 0 81424 400 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 82208 0 82264 400 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 83048 0 83104 400 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 83888 0 83944 400 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 84728 0 84784 400 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 85568 0 85624 400 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 40208 0 40264 400 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 86408 0 86464 400 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 87248 0 87304 400 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 88088 0 88144 400 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 88928 0 88984 400 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 89768 0 89824 400 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 90608 0 90664 400 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 91448 0 91504 400 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 92288 0 92344 400 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 93128 0 93184 400 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 93968 0 94024 400 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 41048 0 41104 400 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 94808 0 94864 400 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 95648 0 95704 400 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 96488 0 96544 400 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 98168 0 98224 400 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 99008 0 99064 400 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 99848 0 99904 400 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 100688 0 100744 400 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 101528 0 101584 400 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 102368 0 102424 400 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 103208 0 103264 400 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 104888 0 104944 400 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 105728 0 105784 400 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 106568 0 106624 400 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 107408 0 107464 400 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 108248 0 108304 400 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 109088 0 109144 400 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 109928 0 109984 400 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 110768 0 110824 400 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 42728 0 42784 400 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 111608 0 111664 400 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 112448 0 112504 400 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 113288 0 113344 400 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 114128 0 114184 400 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 114968 0 115024 400 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 115808 0 115864 400 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 116648 0 116704 400 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 118328 0 118384 400 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 119168 0 119224 400 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 43568 0 43624 400 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 120288 0 120344 400 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 121128 0 121184 400 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 122808 0 122864 400 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 123648 0 123704 400 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 124488 0 124544 400 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 125328 0 125384 400 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 126168 0 126224 400 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 127008 0 127064 400 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 127848 0 127904 400 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 128688 0 128744 400 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 129528 0 129584 400 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 130368 0 130424 400 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 131208 0 131264 400 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 132048 0 132104 400 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 132888 0 132944 400 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 133728 0 133784 400 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 134568 0 134624 400 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 136248 0 136304 400 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 45528 0 45584 400 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 137088 0 137144 400 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 137928 0 137984 400 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 138768 0 138824 400 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 139608 0 139664 400 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 140448 0 140504 400 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 141288 0 141344 400 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 142128 0 142184 400 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 142968 0 143024 400 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 47208 0 47264 400 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 48888 0 48944 400 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 50568 0 50624 400 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 51408 0 51464 400 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 52248 0 52304 400 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 37128 0 37184 400 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 53928 0 53984 400 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 55608 0 55664 400 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 56448 0 56504 400 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 57288 0 57344 400 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 58128 0 58184 400 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 58968 0 59024 400 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 60648 0 60704 400 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 62328 0 62384 400 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 63168 0 63224 400 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 64008 0 64064 400 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 64848 0 64904 400 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 65688 0 65744 400 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 67368 0 67424 400 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 69048 0 69104 400 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 38808 0 38864 400 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 69888 0 69944 400 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 70728 0 70784 400 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 72408 0 72464 400 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 74088 0 74144 400 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 75768 0 75824 400 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 76608 0 76664 400 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 77448 0 77504 400 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 78288 0 78344 400 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 79128 0 79184 400 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 79968 0 80024 400 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 80808 0 80864 400 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 82488 0 82544 400 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 83328 0 83384 400 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 84168 0 84224 400 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 85008 0 85064 400 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 85848 0 85904 400 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 40488 0 40544 400 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 86688 0 86744 400 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 87528 0 87584 400 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 89208 0 89264 400 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 90048 0 90104 400 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 90888 0 90944 400 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 91728 0 91784 400 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 92568 0 92624 400 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 93408 0 93464 400 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 94248 0 94304 400 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 95088 0 95144 400 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 95928 0 95984 400 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 96768 0 96824 400 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 97608 0 97664 400 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 98448 0 98504 400 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 99288 0 99344 400 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 100128 0 100184 400 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 100968 0 101024 400 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 101808 0 101864 400 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 102648 0 102704 400 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 42168 0 42224 400 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 103488 0 103544 400 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 104328 0 104384 400 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 105168 0 105224 400 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 106008 0 106064 400 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 106848 0 106904 400 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 107688 0 107744 400 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 109368 0 109424 400 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 110208 0 110264 400 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 111048 0 111104 400 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 43008 0 43064 400 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 111888 0 111944 400 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 112728 0 112784 400 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 113568 0 113624 400 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 114408 0 114464 400 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 116088 0 116144 400 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 116928 0 116984 400 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 117768 0 117824 400 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 118608 0 118664 400 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 119448 0 119504 400 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 43848 0 43904 400 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 2224 1538 2384 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 6048 0 6104 400 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 6328 0 6384 400 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 18088 0 18144 400 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 19768 0 19824 400 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 20608 0 20664 400 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 21448 0 21504 400 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 23128 0 23184 400 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 24808 0 24864 400 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 26488 0 26544 400 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 28168 0 28224 400 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 29848 0 29904 400 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 31528 0 31584 400 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 33208 0 33264 400 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 13048 0 13104 400 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 14728 0 14784 400 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 15568 0 15624 400 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 16408 0 16464 400 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 17528 0 17584 400 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 19208 0 19264 400 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 20888 0 20944 400 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 22568 0 22624 400 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 24248 0 24304 400 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 9128 0 9184 400 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 25928 0 25984 400 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 27608 0 27664 400 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 29288 0 29344 400 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 30968 0 31024 400 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 32648 0 32704 400 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 10248 0 10304 400 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 34328 0 34384 400 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 11368 0 11424 400 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 12488 0 12544 400 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14168 0 14224 400 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 15848 0 15904 400 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 18648 0 18704 400 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 20328 0 20384 400 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 22008 0 22064 400 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 22848 0 22904 400 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 23688 0 23744 400 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 25368 0 25424 400 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 27048 0 27104 400 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 28728 0 28784 400 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 29568 0 29624 400 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 30408 0 30464 400 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 31248 0 31304 400 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 32088 0 32144 400 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 33768 0 33824 400 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 35448 0 35504 400 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 11648 0 11704 400 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 13608 0 13664 400 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 15288 0 15344 400 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 16968 0 17024 400 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 8568 0 8624 400 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 9688 0 9744 400 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 10808 0 10864 400 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 11928 0 11984 400 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 7448 0 7504 400 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 59928544
string GDS_FILE /home/cra2ypierr0t/workspace/caravel_jacaranda-8_GF180/openlane/computer/runs/22_12_04_19_43/results/signoff/computer.magic.gds
string GDS_START 517410
<< end >>

