VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3000.000 BY 3000.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1216.600 3004.800 1217.720 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2286.760 2997.600 2287.880 3004.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1955.240 2997.600 1956.360 3004.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1623.720 2997.600 1624.840 3004.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1292.200 2997.600 1293.320 3004.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.680 2997.600 961.800 3004.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 629.160 2997.600 630.280 3004.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.640 2997.600 298.760 3004.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2968.280 2.400 2969.400 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2746.520 2.400 2747.640 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2524.760 2.400 2525.880 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1442.840 3004.800 1443.960 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2303.000 2.400 2304.120 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2081.240 2.400 2082.360 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1859.480 2.400 1860.600 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1637.720 2.400 1638.840 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1415.960 2.400 1417.080 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1194.200 2.400 1195.320 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 972.440 2.400 973.560 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 750.680 2.400 751.800 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 528.920 2.400 530.040 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1669.080 3004.800 1670.200 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1895.320 3004.800 1896.440 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2121.560 3004.800 2122.680 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2347.800 3004.800 2348.920 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2574.040 3004.800 2575.160 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2800.280 3004.800 2801.400 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2949.800 2997.600 2950.920 3004.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2618.280 2997.600 2619.400 3004.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 28.840 3004.800 29.960 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1951.880 3004.800 1953.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2178.120 3004.800 2179.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2404.360 3004.800 2405.480 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2630.600 3004.800 2631.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2856.840 3004.800 2857.960 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2866.920 2997.600 2868.040 3004.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2535.400 2997.600 2536.520 3004.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2203.880 2997.600 2205.000 3004.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1872.360 2997.600 1873.480 3004.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1540.840 2997.600 1541.960 3004.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 198.520 3004.800 199.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1209.320 2997.600 1210.440 3004.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 877.800 2997.600 878.920 3004.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.280 2997.600 547.400 3004.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.760 2997.600 215.880 3004.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2912.840 2.400 2913.960 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2691.080 2.400 2692.200 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2469.320 2.400 2470.440 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2247.560 2.400 2248.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2025.800 2.400 2026.920 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1804.040 2.400 1805.160 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 368.200 3004.800 369.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1582.280 2.400 1583.400 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1360.520 2.400 1361.640 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1138.760 2.400 1139.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 917.000 2.400 918.120 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 695.240 2.400 696.360 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 473.480 2.400 474.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 307.160 2.400 308.280 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 140.840 2.400 141.960 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 537.880 3004.800 539.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 707.560 3004.800 708.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 877.240 3004.800 878.360 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1046.920 3004.800 1048.040 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1273.160 3004.800 1274.280 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1499.400 3004.800 1500.520 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1725.640 3004.800 1726.760 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 141.960 3004.800 143.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2065.000 3004.800 2066.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2291.240 3004.800 2292.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2517.480 3004.800 2518.600 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2743.720 3004.800 2744.840 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2969.960 3004.800 2971.080 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2701.160 2997.600 2702.280 3004.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2369.640 2997.600 2370.760 3004.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2038.120 2997.600 2039.240 3004.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1706.600 2997.600 1707.720 3004.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1375.080 2997.600 1376.200 3004.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 311.640 3004.800 312.760 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1043.560 2997.600 1044.680 3004.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.040 2997.600 713.160 3004.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.520 2997.600 381.640 3004.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.000 2997.600 50.120 3004.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2801.960 2.400 2803.080 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2580.200 2.400 2581.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2358.440 2.400 2359.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2136.680 2.400 2137.800 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1914.920 2.400 1916.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1693.160 2.400 1694.280 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 481.320 3004.800 482.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1471.400 2.400 1472.520 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1249.640 2.400 1250.760 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1027.880 2.400 1029.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 806.120 2.400 807.240 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 584.360 2.400 585.480 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 362.600 2.400 363.720 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 196.280 2.400 197.400 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 29.960 2.400 31.080 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 651.000 3004.800 652.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 820.680 3004.800 821.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 990.360 3004.800 991.480 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1160.040 3004.800 1161.160 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1386.280 3004.800 1387.400 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1612.520 3004.800 1613.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1838.760 3004.800 1839.880 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 85.400 3004.800 86.520 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2008.440 3004.800 2009.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2234.680 3004.800 2235.800 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2460.920 3004.800 2462.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2687.160 3004.800 2688.280 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2913.400 3004.800 2914.520 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2784.040 2997.600 2785.160 3004.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2452.520 2997.600 2453.640 3004.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2121.000 2997.600 2122.120 3004.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1789.480 2997.600 1790.600 3004.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1457.960 2997.600 1459.080 3004.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 255.080 3004.800 256.200 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1126.440 2997.600 1127.560 3004.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.920 2997.600 796.040 3004.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.400 2997.600 464.520 3004.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.880 2997.600 133.000 3004.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2857.400 2.400 2858.520 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2635.640 2.400 2636.760 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2413.880 2.400 2415.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2192.120 2.400 2193.240 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1970.360 2.400 1971.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1748.600 2.400 1749.720 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 424.760 3004.800 425.880 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1526.840 2.400 1527.960 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1305.080 2.400 1306.200 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1083.320 2.400 1084.440 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 861.560 2.400 862.680 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 639.800 2.400 640.920 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 418.040 2.400 419.160 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 251.720 2.400 252.840 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 85.400 2.400 86.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 594.440 3004.800 595.560 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 764.120 3004.800 765.240 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 933.800 3004.800 934.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1103.480 3004.800 1104.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1329.720 3004.800 1330.840 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1555.960 3004.800 1557.080 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1782.200 3004.800 1783.320 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.600 -4.800 713.720 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2392.600 -4.800 2393.720 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2409.400 -4.800 2410.520 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2426.200 -4.800 2427.320 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2443.000 -4.800 2444.120 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2459.800 -4.800 2460.920 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2476.600 -4.800 2477.720 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2493.400 -4.800 2494.520 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2510.200 -4.800 2511.320 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2527.000 -4.800 2528.120 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2543.800 -4.800 2544.920 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.600 -4.800 881.720 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2560.600 -4.800 2561.720 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2577.400 -4.800 2578.520 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2594.200 -4.800 2595.320 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2611.000 -4.800 2612.120 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2627.800 -4.800 2628.920 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2644.600 -4.800 2645.720 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2661.400 -4.800 2662.520 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2678.200 -4.800 2679.320 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2695.000 -4.800 2696.120 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2711.800 -4.800 2712.920 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.400 -4.800 898.520 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2728.600 -4.800 2729.720 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2745.400 -4.800 2746.520 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2762.200 -4.800 2763.320 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2779.000 -4.800 2780.120 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2795.800 -4.800 2796.920 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2812.600 -4.800 2813.720 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2829.400 -4.800 2830.520 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2846.200 -4.800 2847.320 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 914.200 -4.800 915.320 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 931.000 -4.800 932.120 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.800 -4.800 948.920 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.600 -4.800 965.720 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.400 -4.800 982.520 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 998.200 -4.800 999.320 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1015.000 -4.800 1016.120 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1031.800 -4.800 1032.920 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.400 -4.800 730.520 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.600 -4.800 1049.720 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.400 -4.800 1066.520 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1082.200 -4.800 1083.320 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1099.000 -4.800 1100.120 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1115.800 -4.800 1116.920 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.600 -4.800 1133.720 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1149.400 -4.800 1150.520 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1166.200 -4.800 1167.320 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1183.000 -4.800 1184.120 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1199.800 -4.800 1200.920 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 746.200 -4.800 747.320 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1216.600 -4.800 1217.720 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1233.400 -4.800 1234.520 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1250.200 -4.800 1251.320 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1267.000 -4.800 1268.120 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1283.800 -4.800 1284.920 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1300.600 -4.800 1301.720 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1317.400 -4.800 1318.520 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1334.200 -4.800 1335.320 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1351.000 -4.800 1352.120 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1367.800 -4.800 1368.920 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.000 -4.800 764.120 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1384.600 -4.800 1385.720 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1401.400 -4.800 1402.520 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1418.200 -4.800 1419.320 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1435.000 -4.800 1436.120 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1451.800 -4.800 1452.920 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1468.600 -4.800 1469.720 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1485.400 -4.800 1486.520 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1502.200 -4.800 1503.320 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1519.000 -4.800 1520.120 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1535.800 -4.800 1536.920 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.800 -4.800 780.920 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1552.600 -4.800 1553.720 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1569.400 -4.800 1570.520 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1586.200 -4.800 1587.320 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1603.000 -4.800 1604.120 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1619.800 -4.800 1620.920 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1636.600 -4.800 1637.720 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1653.400 -4.800 1654.520 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1670.200 -4.800 1671.320 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1687.000 -4.800 1688.120 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1703.800 -4.800 1704.920 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 796.600 -4.800 797.720 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1720.600 -4.800 1721.720 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1737.400 -4.800 1738.520 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1754.200 -4.800 1755.320 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1771.000 -4.800 1772.120 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1787.800 -4.800 1788.920 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1804.600 -4.800 1805.720 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1821.400 -4.800 1822.520 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1838.200 -4.800 1839.320 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1855.000 -4.800 1856.120 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1871.800 -4.800 1872.920 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.400 -4.800 814.520 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1888.600 -4.800 1889.720 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1905.400 -4.800 1906.520 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1922.200 -4.800 1923.320 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1939.000 -4.800 1940.120 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1955.800 -4.800 1956.920 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1972.600 -4.800 1973.720 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1989.400 -4.800 1990.520 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2006.200 -4.800 2007.320 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2023.000 -4.800 2024.120 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2039.800 -4.800 2040.920 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 830.200 -4.800 831.320 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2056.600 -4.800 2057.720 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2073.400 -4.800 2074.520 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2090.200 -4.800 2091.320 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2107.000 -4.800 2108.120 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2123.800 -4.800 2124.920 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2140.600 -4.800 2141.720 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2157.400 -4.800 2158.520 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2174.200 -4.800 2175.320 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2191.000 -4.800 2192.120 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2207.800 -4.800 2208.920 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.000 -4.800 848.120 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2224.600 -4.800 2225.720 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2241.400 -4.800 2242.520 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2258.200 -4.800 2259.320 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2275.000 -4.800 2276.120 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2291.800 -4.800 2292.920 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2308.600 -4.800 2309.720 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2325.400 -4.800 2326.520 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2342.200 -4.800 2343.320 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2359.000 -4.800 2360.120 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2375.800 -4.800 2376.920 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.800 -4.800 864.920 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 718.200 -4.800 719.320 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2398.200 -4.800 2399.320 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2415.000 -4.800 2416.120 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2431.800 -4.800 2432.920 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2448.600 -4.800 2449.720 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2465.400 -4.800 2466.520 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2482.200 -4.800 2483.320 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2499.000 -4.800 2500.120 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2515.800 -4.800 2516.920 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2532.600 -4.800 2533.720 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2549.400 -4.800 2550.520 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 886.200 -4.800 887.320 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2566.200 -4.800 2567.320 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2583.000 -4.800 2584.120 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2599.800 -4.800 2600.920 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2616.600 -4.800 2617.720 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2633.400 -4.800 2634.520 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2650.200 -4.800 2651.320 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2667.000 -4.800 2668.120 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2683.800 -4.800 2684.920 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2700.600 -4.800 2701.720 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2717.400 -4.800 2718.520 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.000 -4.800 904.120 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2734.200 -4.800 2735.320 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2751.000 -4.800 2752.120 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2767.800 -4.800 2768.920 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2784.600 -4.800 2785.720 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2801.400 -4.800 2802.520 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2818.200 -4.800 2819.320 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2835.000 -4.800 2836.120 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2851.800 -4.800 2852.920 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 919.800 -4.800 920.920 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 936.600 -4.800 937.720 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 953.400 -4.800 954.520 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 970.200 -4.800 971.320 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 987.000 -4.800 988.120 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1003.800 -4.800 1004.920 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1020.600 -4.800 1021.720 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.400 -4.800 1038.520 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.000 -4.800 736.120 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1054.200 -4.800 1055.320 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.000 -4.800 1072.120 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1087.800 -4.800 1088.920 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1104.600 -4.800 1105.720 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1121.400 -4.800 1122.520 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1138.200 -4.800 1139.320 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1155.000 -4.800 1156.120 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1171.800 -4.800 1172.920 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1188.600 -4.800 1189.720 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1205.400 -4.800 1206.520 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.800 -4.800 752.920 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1222.200 -4.800 1223.320 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1239.000 -4.800 1240.120 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1255.800 -4.800 1256.920 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1272.600 -4.800 1273.720 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1289.400 -4.800 1290.520 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1306.200 -4.800 1307.320 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1323.000 -4.800 1324.120 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1339.800 -4.800 1340.920 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1356.600 -4.800 1357.720 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1373.400 -4.800 1374.520 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 768.600 -4.800 769.720 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1390.200 -4.800 1391.320 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1407.000 -4.800 1408.120 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1423.800 -4.800 1424.920 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1440.600 -4.800 1441.720 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1457.400 -4.800 1458.520 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1474.200 -4.800 1475.320 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1491.000 -4.800 1492.120 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1507.800 -4.800 1508.920 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1524.600 -4.800 1525.720 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1541.400 -4.800 1542.520 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 785.400 -4.800 786.520 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1558.200 -4.800 1559.320 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1575.000 -4.800 1576.120 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1591.800 -4.800 1592.920 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1608.600 -4.800 1609.720 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1625.400 -4.800 1626.520 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1642.200 -4.800 1643.320 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1659.000 -4.800 1660.120 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1675.800 -4.800 1676.920 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1692.600 -4.800 1693.720 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1709.400 -4.800 1710.520 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 802.200 -4.800 803.320 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1726.200 -4.800 1727.320 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1743.000 -4.800 1744.120 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1759.800 -4.800 1760.920 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1776.600 -4.800 1777.720 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1793.400 -4.800 1794.520 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1810.200 -4.800 1811.320 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1827.000 -4.800 1828.120 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1843.800 -4.800 1844.920 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1860.600 -4.800 1861.720 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1877.400 -4.800 1878.520 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.000 -4.800 820.120 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1894.200 -4.800 1895.320 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1911.000 -4.800 1912.120 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1927.800 -4.800 1928.920 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1944.600 -4.800 1945.720 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1961.400 -4.800 1962.520 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1978.200 -4.800 1979.320 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1995.000 -4.800 1996.120 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2011.800 -4.800 2012.920 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2028.600 -4.800 2029.720 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2045.400 -4.800 2046.520 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 835.800 -4.800 836.920 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2062.200 -4.800 2063.320 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2079.000 -4.800 2080.120 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2095.800 -4.800 2096.920 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2112.600 -4.800 2113.720 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2129.400 -4.800 2130.520 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2146.200 -4.800 2147.320 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2163.000 -4.800 2164.120 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2179.800 -4.800 2180.920 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2196.600 -4.800 2197.720 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2213.400 -4.800 2214.520 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 852.600 -4.800 853.720 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2230.200 -4.800 2231.320 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2247.000 -4.800 2248.120 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2263.800 -4.800 2264.920 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2280.600 -4.800 2281.720 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2297.400 -4.800 2298.520 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2314.200 -4.800 2315.320 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2331.000 -4.800 2332.120 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2347.800 -4.800 2348.920 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2364.600 -4.800 2365.720 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2381.400 -4.800 2382.520 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 869.400 -4.800 870.520 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.800 -4.800 724.920 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2403.800 -4.800 2404.920 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2420.600 -4.800 2421.720 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2437.400 -4.800 2438.520 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2454.200 -4.800 2455.320 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2471.000 -4.800 2472.120 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2487.800 -4.800 2488.920 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2504.600 -4.800 2505.720 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2521.400 -4.800 2522.520 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2538.200 -4.800 2539.320 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2555.000 -4.800 2556.120 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 891.800 -4.800 892.920 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2571.800 -4.800 2572.920 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2588.600 -4.800 2589.720 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2605.400 -4.800 2606.520 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2622.200 -4.800 2623.320 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2639.000 -4.800 2640.120 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2655.800 -4.800 2656.920 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2672.600 -4.800 2673.720 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2689.400 -4.800 2690.520 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2706.200 -4.800 2707.320 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2723.000 -4.800 2724.120 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 908.600 -4.800 909.720 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2739.800 -4.800 2740.920 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2756.600 -4.800 2757.720 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2773.400 -4.800 2774.520 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2790.200 -4.800 2791.320 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2807.000 -4.800 2808.120 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2823.800 -4.800 2824.920 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2840.600 -4.800 2841.720 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2857.400 -4.800 2858.520 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 925.400 -4.800 926.520 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 942.200 -4.800 943.320 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 959.000 -4.800 960.120 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 975.800 -4.800 976.920 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 992.600 -4.800 993.720 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1009.400 -4.800 1010.520 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1026.200 -4.800 1027.320 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1043.000 -4.800 1044.120 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 740.600 -4.800 741.720 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1059.800 -4.800 1060.920 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1076.600 -4.800 1077.720 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1093.400 -4.800 1094.520 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1110.200 -4.800 1111.320 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1127.000 -4.800 1128.120 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1143.800 -4.800 1144.920 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1160.600 -4.800 1161.720 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1177.400 -4.800 1178.520 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1194.200 -4.800 1195.320 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1211.000 -4.800 1212.120 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 757.400 -4.800 758.520 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1227.800 -4.800 1228.920 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1244.600 -4.800 1245.720 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1261.400 -4.800 1262.520 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1278.200 -4.800 1279.320 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1295.000 -4.800 1296.120 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1311.800 -4.800 1312.920 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1328.600 -4.800 1329.720 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1345.400 -4.800 1346.520 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1362.200 -4.800 1363.320 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1379.000 -4.800 1380.120 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 774.200 -4.800 775.320 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1395.800 -4.800 1396.920 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1412.600 -4.800 1413.720 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1429.400 -4.800 1430.520 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1446.200 -4.800 1447.320 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1463.000 -4.800 1464.120 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1479.800 -4.800 1480.920 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1496.600 -4.800 1497.720 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1513.400 -4.800 1514.520 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1530.200 -4.800 1531.320 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1547.000 -4.800 1548.120 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 791.000 -4.800 792.120 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1563.800 -4.800 1564.920 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1580.600 -4.800 1581.720 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1597.400 -4.800 1598.520 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1614.200 -4.800 1615.320 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1631.000 -4.800 1632.120 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1647.800 -4.800 1648.920 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1664.600 -4.800 1665.720 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1681.400 -4.800 1682.520 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1698.200 -4.800 1699.320 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1715.000 -4.800 1716.120 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 807.800 -4.800 808.920 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1731.800 -4.800 1732.920 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1748.600 -4.800 1749.720 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1765.400 -4.800 1766.520 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1782.200 -4.800 1783.320 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1799.000 -4.800 1800.120 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1815.800 -4.800 1816.920 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1832.600 -4.800 1833.720 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1849.400 -4.800 1850.520 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1866.200 -4.800 1867.320 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1883.000 -4.800 1884.120 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 824.600 -4.800 825.720 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1899.800 -4.800 1900.920 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1916.600 -4.800 1917.720 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1933.400 -4.800 1934.520 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1950.200 -4.800 1951.320 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1967.000 -4.800 1968.120 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1983.800 -4.800 1984.920 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2000.600 -4.800 2001.720 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2017.400 -4.800 2018.520 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2034.200 -4.800 2035.320 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2051.000 -4.800 2052.120 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 841.400 -4.800 842.520 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2067.800 -4.800 2068.920 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2084.600 -4.800 2085.720 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2101.400 -4.800 2102.520 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2118.200 -4.800 2119.320 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2135.000 -4.800 2136.120 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2151.800 -4.800 2152.920 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2168.600 -4.800 2169.720 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2185.400 -4.800 2186.520 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2202.200 -4.800 2203.320 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2219.000 -4.800 2220.120 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 858.200 -4.800 859.320 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2235.800 -4.800 2236.920 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2252.600 -4.800 2253.720 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2269.400 -4.800 2270.520 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2286.200 -4.800 2287.320 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2303.000 -4.800 2304.120 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2319.800 -4.800 2320.920 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2336.600 -4.800 2337.720 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2353.400 -4.800 2354.520 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.200 -4.800 2371.320 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2387.000 -4.800 2388.120 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.000 -4.800 876.120 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2863.000 -4.800 2864.120 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2868.600 -4.800 2869.720 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2874.200 -4.800 2875.320 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2879.800 -4.800 2880.920 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -8.830 0.130 -5.730 2998.670 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -8.830 0.130 3008.750 3.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -8.830 2995.570 3008.750 2998.670 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3005.650 0.130 3008.750 2998.670 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 10.170 -33.470 13.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.170 -33.470 193.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.170 -33.470 373.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.170 -33.470 553.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 730.170 -33.470 733.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 730.170 2335.270 733.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 910.170 -33.470 913.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 910.170 2335.270 913.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1090.170 -33.470 1093.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1090.170 2335.270 1093.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1270.170 -33.470 1273.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1270.170 2335.270 1273.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1450.170 -33.470 1453.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1450.170 2335.270 1453.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1630.170 -33.470 1633.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1630.170 2335.270 1633.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1810.170 -33.470 1813.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1810.170 2335.270 1813.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1990.170 -33.470 1993.270 850.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1990.170 2337.340 1993.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.170 -33.470 2173.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2350.170 -33.470 2353.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2530.170 -33.470 2533.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.170 -33.470 2713.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2890.170 -33.470 2893.270 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 19.130 3042.350 22.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 199.130 3042.350 202.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 379.130 3042.350 382.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 559.130 3042.350 562.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 739.130 3042.350 742.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 919.130 3042.350 922.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1099.130 597.820 1102.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1279.130 597.820 1282.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1459.130 597.820 1462.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1639.130 597.820 1642.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1819.130 597.820 1822.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1999.130 597.820 2002.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2179.130 597.820 2182.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2359.130 3042.350 2362.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2539.130 3042.350 2542.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2719.130 3042.350 2722.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2899.130 3042.350 2902.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1099.130 3042.350 1102.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1279.130 3042.350 1282.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1459.130 3042.350 1462.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1639.130 3042.350 1642.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1819.130 3042.350 1822.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1999.130 3042.350 2002.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2179.130 3042.350 2182.230 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -18.430 -9.470 -15.330 3008.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -18.430 -9.470 3018.350 -6.370 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -18.430 3005.170 3018.350 3008.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3015.250 -9.470 3018.350 3008.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 47.370 -33.470 50.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 227.370 -33.470 230.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 407.370 -33.470 410.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 587.370 -33.470 590.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 767.370 -33.470 770.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 767.370 2335.270 770.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 947.370 -33.470 950.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 947.370 2335.270 950.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.370 -33.470 1130.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.370 2335.270 1130.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1307.370 -33.470 1310.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1307.370 2335.270 1310.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1487.370 -33.470 1490.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1487.370 2335.270 1490.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1667.370 -33.470 1670.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1667.370 2335.270 1670.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1847.370 -33.470 1850.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1847.370 2335.270 1850.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2027.370 -33.470 2030.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2207.370 -33.470 2210.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2387.370 -33.470 2390.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2567.370 -33.470 2570.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2747.370 -33.470 2750.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2927.370 -33.470 2930.470 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 56.330 3042.350 59.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 236.330 3042.350 239.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 416.330 3042.350 419.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 596.330 3042.350 599.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 776.330 3042.350 779.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 956.330 3042.350 959.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1136.330 597.820 1139.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1316.330 597.820 1319.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1496.330 597.820 1499.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1676.330 597.820 1679.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1856.330 597.820 1859.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2036.330 597.820 2039.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2216.330 597.820 2219.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2396.330 3042.350 2399.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2576.330 3042.350 2579.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2756.330 3042.350 2759.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2936.330 3042.350 2939.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1136.330 3042.350 1139.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1316.330 3042.350 1319.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1496.330 3042.350 1499.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1676.330 3042.350 1679.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1856.330 3042.350 1859.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2036.330 3042.350 2039.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2216.330 3042.350 2219.430 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -28.030 -19.070 -24.930 3017.870 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -28.030 -19.070 3027.950 -15.970 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -28.030 3014.770 3027.950 3017.870 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3024.850 -19.070 3027.950 3017.870 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 84.570 -33.470 87.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 264.570 -33.470 267.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 444.570 -33.470 447.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 624.570 -33.470 627.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 624.570 2335.270 627.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 804.570 -33.470 807.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 804.570 2335.270 807.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 984.570 -33.470 987.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 984.570 2335.270 987.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1164.570 -33.470 1167.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1164.570 2335.270 1167.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1344.570 -33.470 1347.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1344.570 2335.270 1347.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1524.570 -33.470 1527.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1524.570 2335.270 1527.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.570 -33.470 1707.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1704.570 2335.270 1707.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1884.570 -33.470 1887.670 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1884.570 2335.270 1887.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2064.570 -33.470 2067.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2244.570 -33.470 2247.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2424.570 -33.470 2427.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2604.570 -33.470 2607.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2784.570 -33.470 2787.670 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2964.570 -33.470 2967.670 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 93.530 3042.350 96.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 273.530 3042.350 276.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 453.530 3042.350 456.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 633.530 3042.350 636.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 813.530 3042.350 816.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 993.530 3042.350 996.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1173.530 597.820 1176.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1353.530 597.820 1356.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1533.530 597.820 1536.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1713.530 597.820 1716.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1893.530 597.820 1896.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2073.530 597.820 2076.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2253.530 597.820 2256.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2433.530 3042.350 2436.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2613.530 3042.350 2616.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2793.530 3042.350 2796.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2973.530 3042.350 2976.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1173.530 3042.350 1176.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1353.530 3042.350 1356.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1533.530 3042.350 1536.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1713.530 3042.350 1716.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1893.530 3042.350 1896.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2073.530 3042.350 2076.630 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2253.530 3042.350 2256.630 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -37.630 -28.670 -34.530 3027.470 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -37.630 -28.670 3037.550 -25.570 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -37.630 3024.370 3037.550 3027.470 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3034.450 -28.670 3037.550 3027.470 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.770 -33.470 124.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 301.770 -33.470 304.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 481.770 -33.470 484.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 661.770 -33.470 664.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 661.770 2335.270 664.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 841.770 -33.470 844.870 850.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 841.770 2337.340 844.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1021.770 -33.470 1024.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1021.770 2335.270 1024.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1201.770 -33.470 1204.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1201.770 2335.270 1204.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1381.770 -33.470 1384.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1381.770 2335.270 1384.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1561.770 -33.470 1564.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1561.770 2335.270 1564.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1741.770 -33.470 1744.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1741.770 2335.270 1744.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1921.770 -33.470 1924.870 851.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1921.770 2335.270 1924.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2101.770 -33.470 2104.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2281.770 -33.470 2284.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2461.770 -33.470 2464.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2641.770 -33.470 2644.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2821.770 -33.470 2824.870 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 130.730 3042.350 133.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 310.730 3042.350 313.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 490.730 3042.350 493.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 670.730 3042.350 673.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 850.730 3042.350 853.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1030.730 597.820 1033.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1210.730 597.820 1213.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1390.730 597.820 1393.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1570.730 597.820 1573.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1750.730 597.820 1753.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1930.730 597.820 1933.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2110.730 597.820 2113.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2290.730 597.820 2293.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2470.730 3042.350 2473.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2650.730 3042.350 2653.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2830.730 3042.350 2833.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1030.730 3042.350 1033.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1210.730 3042.350 1213.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1390.730 3042.350 1393.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1570.730 3042.350 1573.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1750.730 3042.350 1753.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1930.730 3042.350 1933.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2110.730 3042.350 2113.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2290.730 3042.350 2293.830 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -32.830 -23.870 -29.730 3022.670 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -32.830 -23.870 3032.750 -20.770 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -32.830 3019.570 3032.750 3022.670 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3029.650 -23.870 3032.750 3022.670 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.170 -33.470 106.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 283.170 -33.470 286.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 463.170 -33.470 466.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 643.170 -33.470 646.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 643.170 2335.270 646.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 823.170 -33.470 826.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 823.170 2335.270 826.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1003.170 -33.470 1006.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1003.170 2335.270 1006.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1183.170 -33.470 1186.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1183.170 2335.270 1186.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1363.170 -33.470 1366.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1363.170 2335.270 1366.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1543.170 -33.470 1546.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1543.170 2335.270 1546.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1723.170 -33.470 1726.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1723.170 2335.270 1726.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1903.170 -33.470 1906.270 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1903.170 2335.270 1906.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2083.170 -33.470 2086.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2263.170 -33.470 2266.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2443.170 -33.470 2446.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2623.170 -33.470 2626.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2803.170 -33.470 2806.270 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2983.170 -33.470 2986.270 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 112.130 3042.350 115.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 292.130 3042.350 295.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 472.130 3042.350 475.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 652.130 3042.350 655.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 832.130 3042.350 835.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1012.130 597.820 1015.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1192.130 597.820 1195.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1372.130 597.820 1375.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1552.130 597.820 1555.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1732.130 597.820 1735.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1912.130 597.820 1915.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2092.130 597.820 2095.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2272.130 597.820 2275.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2452.130 3042.350 2455.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2632.130 3042.350 2635.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2812.130 3042.350 2815.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1012.130 3042.350 1015.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1192.130 3042.350 1195.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1372.130 3042.350 1375.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1552.130 3042.350 1555.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1732.130 3042.350 1735.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1912.130 3042.350 1915.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2092.130 3042.350 2095.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2272.130 3042.350 2275.230 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -42.430 -33.470 -39.330 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 -33.470 3042.350 -30.370 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 3029.170 3042.350 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3039.250 -33.470 3042.350 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 140.370 -33.470 143.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 320.370 -33.470 323.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 500.370 -33.470 503.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 680.370 -33.470 683.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 680.370 2335.270 683.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 860.370 -33.470 863.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 860.370 2335.270 863.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1040.370 -33.470 1043.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1040.370 2335.270 1043.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1220.370 -33.470 1223.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1220.370 2335.270 1223.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1400.370 -33.470 1403.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1400.370 2335.270 1403.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1580.370 -33.470 1583.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1580.370 2335.270 1583.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1760.370 -33.470 1763.470 850.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1760.370 2337.340 1763.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1940.370 -33.470 1943.470 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1940.370 2335.270 1943.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2120.370 -33.470 2123.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2300.370 -33.470 2303.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2480.370 -33.470 2483.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2660.370 -33.470 2663.470 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2840.370 -33.470 2843.470 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 149.330 3042.350 152.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 329.330 3042.350 332.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 509.330 3042.350 512.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 689.330 3042.350 692.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 869.330 3042.350 872.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1049.330 597.820 1052.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1229.330 597.820 1232.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1409.330 597.820 1412.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1589.330 597.820 1592.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1769.330 597.820 1772.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1949.330 597.820 1952.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2129.330 597.820 2132.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2309.330 3042.350 2312.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2489.330 3042.350 2492.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2669.330 3042.350 2672.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2849.330 3042.350 2852.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1049.330 3042.350 1052.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1229.330 3042.350 1232.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1409.330 3042.350 1412.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1589.330 3042.350 1592.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1769.330 3042.350 1772.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1949.330 3042.350 1952.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2129.330 3042.350 2132.430 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -13.630 -4.670 -10.530 3003.470 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -13.630 -4.670 3013.550 -1.570 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -13.630 3000.370 3013.550 3003.470 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3010.450 -4.670 3013.550 3003.470 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.770 -33.470 31.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.770 -33.470 211.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 388.770 -33.470 391.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.770 -33.470 571.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 748.770 -33.470 751.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 748.770 2335.270 751.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.770 -33.470 931.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.770 2335.270 931.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1108.770 -33.470 1111.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1108.770 2335.270 1111.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1288.770 -33.470 1291.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1288.770 2335.270 1291.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1468.770 -33.470 1471.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1468.770 2335.270 1471.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.770 -33.470 1651.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.770 2335.270 1651.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1828.770 -33.470 1831.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1828.770 2335.270 1831.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2008.770 -33.470 2011.870 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2008.770 2335.270 2011.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2188.770 -33.470 2191.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.770 -33.470 2371.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2548.770 -33.470 2551.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2728.770 -33.470 2731.870 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2908.770 -33.470 2911.870 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 37.730 3042.350 40.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 217.730 3042.350 220.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 397.730 3042.350 400.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 577.730 3042.350 580.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 757.730 3042.350 760.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 937.730 3042.350 940.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1117.730 597.820 1120.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1297.730 597.820 1300.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1477.730 597.820 1480.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1657.730 597.820 1660.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1837.730 597.820 1840.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2017.730 597.820 2020.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2197.730 597.820 2200.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2377.730 3042.350 2380.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2557.730 3042.350 2560.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2737.730 3042.350 2740.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2917.730 3042.350 2920.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1117.730 3042.350 1120.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1297.730 3042.350 1300.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1477.730 3042.350 1480.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1657.730 3042.350 1660.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1837.730 3042.350 1840.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2017.730 3042.350 2020.830 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2197.730 3042.350 2200.830 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -23.230 -14.270 -20.130 3013.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -23.230 -14.270 3023.150 -11.170 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -23.230 3009.970 3023.150 3013.070 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3020.050 -14.270 3023.150 3013.070 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 65.970 -33.470 69.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 245.970 -33.470 249.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 425.970 -33.470 429.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.970 -33.470 609.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.970 2335.270 609.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.970 -33.470 789.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 785.970 2335.270 789.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 965.970 -33.470 969.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 965.970 2335.270 969.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1145.970 -33.470 1149.070 850.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1145.970 2337.340 1149.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1325.970 -33.470 1329.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1325.970 2335.270 1329.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1505.970 -33.470 1509.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1505.970 2335.270 1509.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1685.970 -33.470 1689.070 850.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1685.970 2337.340 1689.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.970 -33.470 1869.070 851.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.970 2335.270 1869.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2045.970 -33.470 2049.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2225.970 -33.470 2229.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2405.970 -33.470 2409.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2585.970 -33.470 2589.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2765.970 -33.470 2769.070 3032.270 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2945.970 -33.470 2949.070 3032.270 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 74.930 3042.350 78.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 254.930 3042.350 258.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 434.930 3042.350 438.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 614.930 3042.350 618.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 794.930 3042.350 798.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 974.930 3042.350 978.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1154.930 597.820 1158.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1334.930 597.820 1338.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1514.930 597.820 1518.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1694.930 597.820 1698.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 1874.930 597.820 1878.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2054.930 597.820 2058.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2234.930 597.820 2238.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2414.930 3042.350 2418.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2594.930 3042.350 2598.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2774.930 3042.350 2778.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -42.430 2954.930 3042.350 2958.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1154.930 3042.350 1158.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1334.930 3042.350 1338.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1514.930 3042.350 1518.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1694.930 3042.350 1698.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 1874.930 3042.350 1878.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2054.930 3042.350 2058.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1996.780 2234.930 3042.350 2238.030 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.000 -4.800 120.120 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.600 -4.800 125.720 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 -4.800 131.320 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.600 -4.800 153.720 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.000 -4.800 344.120 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.800 -4.800 360.920 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.600 -4.800 377.720 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.400 -4.800 394.520 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 410.200 -4.800 411.320 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.000 -4.800 428.120 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.800 -4.800 444.920 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.600 -4.800 461.720 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.400 -4.800 478.520 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.200 -4.800 495.320 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.000 -4.800 176.120 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.000 -4.800 512.120 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.800 -4.800 528.920 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.600 -4.800 545.720 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.400 -4.800 562.520 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 578.200 -4.800 579.320 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 595.000 -4.800 596.120 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.800 -4.800 612.920 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.600 -4.800 629.720 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.400 -4.800 646.520 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 662.200 -4.800 663.320 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.400 -4.800 198.520 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 679.000 -4.800 680.120 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 695.800 -4.800 696.920 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.800 -4.800 220.920 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.200 -4.800 243.320 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.000 -4.800 260.120 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 -4.800 276.920 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.600 -4.800 293.720 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.400 -4.800 310.520 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 326.200 -4.800 327.320 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.800 -4.800 136.920 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.200 -4.800 159.320 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.600 -4.800 349.720 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.400 -4.800 366.520 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.200 -4.800 383.320 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.000 -4.800 400.120 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 415.800 -4.800 416.920 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 432.600 -4.800 433.720 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.400 -4.800 450.520 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.200 -4.800 467.320 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.000 -4.800 484.120 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.800 -4.800 500.920 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 -4.800 181.720 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.600 -4.800 517.720 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 533.400 -4.800 534.520 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 550.200 -4.800 551.320 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.000 -4.800 568.120 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 583.800 -4.800 584.920 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 600.600 -4.800 601.720 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 617.400 -4.800 618.520 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 634.200 -4.800 635.320 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.000 -4.800 652.120 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 667.800 -4.800 668.920 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.000 -4.800 204.120 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 684.600 -4.800 685.720 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 701.400 -4.800 702.520 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.400 -4.800 226.520 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.800 -4.800 248.920 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.600 -4.800 265.720 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.400 -4.800 282.520 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.200 -4.800 299.320 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.000 -4.800 316.120 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 331.800 -4.800 332.920 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.800 -4.800 164.920 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 354.200 -4.800 355.320 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 -4.800 372.120 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.800 -4.800 388.920 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 404.600 -4.800 405.720 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.400 -4.800 422.520 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 438.200 -4.800 439.320 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.000 -4.800 456.120 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 471.800 -4.800 472.920 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.600 -4.800 489.720 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.400 -4.800 506.520 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.200 -4.800 187.320 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 522.200 -4.800 523.320 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.000 -4.800 540.120 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 555.800 -4.800 556.920 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.600 -4.800 573.720 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 589.400 -4.800 590.520 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 606.200 -4.800 607.320 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 623.000 -4.800 624.120 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 639.800 -4.800 640.920 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 656.600 -4.800 657.720 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.400 -4.800 674.520 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.600 -4.800 209.720 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 690.200 -4.800 691.320 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 707.000 -4.800 708.120 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.000 -4.800 232.120 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.400 -4.800 254.520 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.200 -4.800 271.320 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.000 -4.800 288.120 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 303.800 -4.800 304.920 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.600 -4.800 321.720 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.400 -4.800 338.520 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.400 -4.800 170.520 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.800 -4.800 192.920 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.200 -4.800 215.320 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.600 -4.800 237.720 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.400 -4.800 142.520 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.000 -4.800 148.120 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 151.290 20.870 2759.030 2327.730 ;
      LAYER Metal2 ;
        RECT 20.300 2997.300 48.700 2998.100 ;
        RECT 50.420 2997.300 131.580 2998.100 ;
        RECT 133.300 2997.300 214.460 2998.100 ;
        RECT 216.180 2997.300 297.340 2998.100 ;
        RECT 299.060 2997.300 380.220 2998.100 ;
        RECT 381.940 2997.300 463.100 2998.100 ;
        RECT 464.820 2997.300 545.980 2998.100 ;
        RECT 547.700 2997.300 628.860 2998.100 ;
        RECT 630.580 2997.300 711.740 2998.100 ;
        RECT 713.460 2997.300 794.620 2998.100 ;
        RECT 796.340 2997.300 877.500 2998.100 ;
        RECT 879.220 2997.300 960.380 2998.100 ;
        RECT 962.100 2997.300 1043.260 2998.100 ;
        RECT 1044.980 2997.300 1126.140 2998.100 ;
        RECT 1127.860 2997.300 1209.020 2998.100 ;
        RECT 1210.740 2997.300 1291.900 2998.100 ;
        RECT 1293.620 2997.300 1374.780 2998.100 ;
        RECT 1376.500 2997.300 1457.660 2998.100 ;
        RECT 1459.380 2997.300 1540.540 2998.100 ;
        RECT 1542.260 2997.300 1623.420 2998.100 ;
        RECT 1625.140 2997.300 1706.300 2998.100 ;
        RECT 1708.020 2997.300 1789.180 2998.100 ;
        RECT 1790.900 2997.300 1872.060 2998.100 ;
        RECT 1873.780 2997.300 1954.940 2998.100 ;
        RECT 1956.660 2997.300 2037.820 2998.100 ;
        RECT 2039.540 2997.300 2120.700 2998.100 ;
        RECT 2122.420 2997.300 2203.580 2998.100 ;
        RECT 2205.300 2997.300 2286.460 2998.100 ;
        RECT 2288.180 2997.300 2369.340 2998.100 ;
        RECT 2371.060 2997.300 2452.220 2998.100 ;
        RECT 2453.940 2997.300 2535.100 2998.100 ;
        RECT 2536.820 2997.300 2617.980 2998.100 ;
        RECT 2619.700 2997.300 2700.860 2998.100 ;
        RECT 2702.580 2997.300 2783.740 2998.100 ;
        RECT 2785.460 2997.300 2866.620 2998.100 ;
        RECT 2868.340 2997.300 2949.500 2998.100 ;
        RECT 2951.220 2997.300 2980.740 2998.100 ;
        RECT 20.300 2.700 2980.740 2997.300 ;
        RECT 20.300 0.090 118.700 2.700 ;
        RECT 120.420 0.090 124.300 2.700 ;
        RECT 126.020 0.090 129.900 2.700 ;
        RECT 131.620 0.090 135.500 2.700 ;
        RECT 137.220 0.090 141.100 2.700 ;
        RECT 142.820 0.090 146.700 2.700 ;
        RECT 148.420 0.090 152.300 2.700 ;
        RECT 154.020 0.090 157.900 2.700 ;
        RECT 159.620 0.090 163.500 2.700 ;
        RECT 165.220 0.090 169.100 2.700 ;
        RECT 170.820 0.090 174.700 2.700 ;
        RECT 176.420 0.090 180.300 2.700 ;
        RECT 182.020 0.090 185.900 2.700 ;
        RECT 187.620 0.090 191.500 2.700 ;
        RECT 193.220 0.090 197.100 2.700 ;
        RECT 198.820 0.090 202.700 2.700 ;
        RECT 204.420 0.090 208.300 2.700 ;
        RECT 210.020 0.090 213.900 2.700 ;
        RECT 215.620 0.090 219.500 2.700 ;
        RECT 221.220 0.090 225.100 2.700 ;
        RECT 226.820 0.090 230.700 2.700 ;
        RECT 232.420 0.090 236.300 2.700 ;
        RECT 238.020 0.090 241.900 2.700 ;
        RECT 243.620 0.090 247.500 2.700 ;
        RECT 249.220 0.090 253.100 2.700 ;
        RECT 254.820 0.090 258.700 2.700 ;
        RECT 260.420 0.090 264.300 2.700 ;
        RECT 266.020 0.090 269.900 2.700 ;
        RECT 271.620 0.090 275.500 2.700 ;
        RECT 277.220 0.090 281.100 2.700 ;
        RECT 282.820 0.090 286.700 2.700 ;
        RECT 288.420 0.090 292.300 2.700 ;
        RECT 294.020 0.090 297.900 2.700 ;
        RECT 299.620 0.090 303.500 2.700 ;
        RECT 305.220 0.090 309.100 2.700 ;
        RECT 310.820 0.090 314.700 2.700 ;
        RECT 316.420 0.090 320.300 2.700 ;
        RECT 322.020 0.090 325.900 2.700 ;
        RECT 327.620 0.090 331.500 2.700 ;
        RECT 333.220 0.090 337.100 2.700 ;
        RECT 338.820 0.090 342.700 2.700 ;
        RECT 344.420 0.090 348.300 2.700 ;
        RECT 350.020 0.090 353.900 2.700 ;
        RECT 355.620 0.090 359.500 2.700 ;
        RECT 361.220 0.090 365.100 2.700 ;
        RECT 366.820 0.090 370.700 2.700 ;
        RECT 372.420 0.090 376.300 2.700 ;
        RECT 378.020 0.090 381.900 2.700 ;
        RECT 383.620 0.090 387.500 2.700 ;
        RECT 389.220 0.090 393.100 2.700 ;
        RECT 394.820 0.090 398.700 2.700 ;
        RECT 400.420 0.090 404.300 2.700 ;
        RECT 406.020 0.090 409.900 2.700 ;
        RECT 411.620 0.090 415.500 2.700 ;
        RECT 417.220 0.090 421.100 2.700 ;
        RECT 422.820 0.090 426.700 2.700 ;
        RECT 428.420 0.090 432.300 2.700 ;
        RECT 434.020 0.090 437.900 2.700 ;
        RECT 439.620 0.090 443.500 2.700 ;
        RECT 445.220 0.090 449.100 2.700 ;
        RECT 450.820 0.090 454.700 2.700 ;
        RECT 456.420 0.090 460.300 2.700 ;
        RECT 462.020 0.090 465.900 2.700 ;
        RECT 467.620 0.090 471.500 2.700 ;
        RECT 473.220 0.090 477.100 2.700 ;
        RECT 478.820 0.090 482.700 2.700 ;
        RECT 484.420 0.090 488.300 2.700 ;
        RECT 490.020 0.090 493.900 2.700 ;
        RECT 495.620 0.090 499.500 2.700 ;
        RECT 501.220 0.090 505.100 2.700 ;
        RECT 506.820 0.090 510.700 2.700 ;
        RECT 512.420 0.090 516.300 2.700 ;
        RECT 518.020 0.090 521.900 2.700 ;
        RECT 523.620 0.090 527.500 2.700 ;
        RECT 529.220 0.090 533.100 2.700 ;
        RECT 534.820 0.090 538.700 2.700 ;
        RECT 540.420 0.090 544.300 2.700 ;
        RECT 546.020 0.090 549.900 2.700 ;
        RECT 551.620 0.090 555.500 2.700 ;
        RECT 557.220 0.090 561.100 2.700 ;
        RECT 562.820 0.090 566.700 2.700 ;
        RECT 568.420 0.090 572.300 2.700 ;
        RECT 574.020 0.090 577.900 2.700 ;
        RECT 579.620 0.090 583.500 2.700 ;
        RECT 585.220 0.090 589.100 2.700 ;
        RECT 590.820 0.090 594.700 2.700 ;
        RECT 596.420 0.090 600.300 2.700 ;
        RECT 602.020 0.090 605.900 2.700 ;
        RECT 607.620 0.090 611.500 2.700 ;
        RECT 613.220 0.090 617.100 2.700 ;
        RECT 618.820 0.090 622.700 2.700 ;
        RECT 624.420 0.090 628.300 2.700 ;
        RECT 630.020 0.090 633.900 2.700 ;
        RECT 635.620 0.090 639.500 2.700 ;
        RECT 641.220 0.090 645.100 2.700 ;
        RECT 646.820 0.090 650.700 2.700 ;
        RECT 652.420 0.090 656.300 2.700 ;
        RECT 658.020 0.090 661.900 2.700 ;
        RECT 663.620 0.090 667.500 2.700 ;
        RECT 669.220 0.090 673.100 2.700 ;
        RECT 674.820 0.090 678.700 2.700 ;
        RECT 680.420 0.090 684.300 2.700 ;
        RECT 686.020 0.090 689.900 2.700 ;
        RECT 691.620 0.090 695.500 2.700 ;
        RECT 697.220 0.090 701.100 2.700 ;
        RECT 702.820 0.090 706.700 2.700 ;
        RECT 708.420 0.090 712.300 2.700 ;
        RECT 714.020 0.090 717.900 2.700 ;
        RECT 719.620 0.090 723.500 2.700 ;
        RECT 725.220 0.090 729.100 2.700 ;
        RECT 730.820 0.090 734.700 2.700 ;
        RECT 736.420 0.090 740.300 2.700 ;
        RECT 742.020 0.090 745.900 2.700 ;
        RECT 747.620 0.090 751.500 2.700 ;
        RECT 753.220 0.090 757.100 2.700 ;
        RECT 758.820 0.090 762.700 2.700 ;
        RECT 764.420 0.090 768.300 2.700 ;
        RECT 770.020 0.090 773.900 2.700 ;
        RECT 775.620 0.090 779.500 2.700 ;
        RECT 781.220 0.090 785.100 2.700 ;
        RECT 786.820 0.090 790.700 2.700 ;
        RECT 792.420 0.090 796.300 2.700 ;
        RECT 798.020 0.090 801.900 2.700 ;
        RECT 803.620 0.090 807.500 2.700 ;
        RECT 809.220 0.090 813.100 2.700 ;
        RECT 814.820 0.090 818.700 2.700 ;
        RECT 820.420 0.090 824.300 2.700 ;
        RECT 826.020 0.090 829.900 2.700 ;
        RECT 831.620 0.090 835.500 2.700 ;
        RECT 837.220 0.090 841.100 2.700 ;
        RECT 842.820 0.090 846.700 2.700 ;
        RECT 848.420 0.090 852.300 2.700 ;
        RECT 854.020 0.090 857.900 2.700 ;
        RECT 859.620 0.090 863.500 2.700 ;
        RECT 865.220 0.090 869.100 2.700 ;
        RECT 870.820 0.090 874.700 2.700 ;
        RECT 876.420 0.090 880.300 2.700 ;
        RECT 882.020 0.090 885.900 2.700 ;
        RECT 887.620 0.090 891.500 2.700 ;
        RECT 893.220 0.090 897.100 2.700 ;
        RECT 898.820 0.090 902.700 2.700 ;
        RECT 904.420 0.090 908.300 2.700 ;
        RECT 910.020 0.090 913.900 2.700 ;
        RECT 915.620 0.090 919.500 2.700 ;
        RECT 921.220 0.090 925.100 2.700 ;
        RECT 926.820 0.090 930.700 2.700 ;
        RECT 932.420 0.090 936.300 2.700 ;
        RECT 938.020 0.090 941.900 2.700 ;
        RECT 943.620 0.090 947.500 2.700 ;
        RECT 949.220 0.090 953.100 2.700 ;
        RECT 954.820 0.090 958.700 2.700 ;
        RECT 960.420 0.090 964.300 2.700 ;
        RECT 966.020 0.090 969.900 2.700 ;
        RECT 971.620 0.090 975.500 2.700 ;
        RECT 977.220 0.090 981.100 2.700 ;
        RECT 982.820 0.090 986.700 2.700 ;
        RECT 988.420 0.090 992.300 2.700 ;
        RECT 994.020 0.090 997.900 2.700 ;
        RECT 999.620 0.090 1003.500 2.700 ;
        RECT 1005.220 0.090 1009.100 2.700 ;
        RECT 1010.820 0.090 1014.700 2.700 ;
        RECT 1016.420 0.090 1020.300 2.700 ;
        RECT 1022.020 0.090 1025.900 2.700 ;
        RECT 1027.620 0.090 1031.500 2.700 ;
        RECT 1033.220 0.090 1037.100 2.700 ;
        RECT 1038.820 0.090 1042.700 2.700 ;
        RECT 1044.420 0.090 1048.300 2.700 ;
        RECT 1050.020 0.090 1053.900 2.700 ;
        RECT 1055.620 0.090 1059.500 2.700 ;
        RECT 1061.220 0.090 1065.100 2.700 ;
        RECT 1066.820 0.090 1070.700 2.700 ;
        RECT 1072.420 0.090 1076.300 2.700 ;
        RECT 1078.020 0.090 1081.900 2.700 ;
        RECT 1083.620 0.090 1087.500 2.700 ;
        RECT 1089.220 0.090 1093.100 2.700 ;
        RECT 1094.820 0.090 1098.700 2.700 ;
        RECT 1100.420 0.090 1104.300 2.700 ;
        RECT 1106.020 0.090 1109.900 2.700 ;
        RECT 1111.620 0.090 1115.500 2.700 ;
        RECT 1117.220 0.090 1121.100 2.700 ;
        RECT 1122.820 0.090 1126.700 2.700 ;
        RECT 1128.420 0.090 1132.300 2.700 ;
        RECT 1134.020 0.090 1137.900 2.700 ;
        RECT 1139.620 0.090 1143.500 2.700 ;
        RECT 1145.220 0.090 1149.100 2.700 ;
        RECT 1150.820 0.090 1154.700 2.700 ;
        RECT 1156.420 0.090 1160.300 2.700 ;
        RECT 1162.020 0.090 1165.900 2.700 ;
        RECT 1167.620 0.090 1171.500 2.700 ;
        RECT 1173.220 0.090 1177.100 2.700 ;
        RECT 1178.820 0.090 1182.700 2.700 ;
        RECT 1184.420 0.090 1188.300 2.700 ;
        RECT 1190.020 0.090 1193.900 2.700 ;
        RECT 1195.620 0.090 1199.500 2.700 ;
        RECT 1201.220 0.090 1205.100 2.700 ;
        RECT 1206.820 0.090 1210.700 2.700 ;
        RECT 1212.420 0.090 1216.300 2.700 ;
        RECT 1218.020 0.090 1221.900 2.700 ;
        RECT 1223.620 0.090 1227.500 2.700 ;
        RECT 1229.220 0.090 1233.100 2.700 ;
        RECT 1234.820 0.090 1238.700 2.700 ;
        RECT 1240.420 0.090 1244.300 2.700 ;
        RECT 1246.020 0.090 1249.900 2.700 ;
        RECT 1251.620 0.090 1255.500 2.700 ;
        RECT 1257.220 0.090 1261.100 2.700 ;
        RECT 1262.820 0.090 1266.700 2.700 ;
        RECT 1268.420 0.090 1272.300 2.700 ;
        RECT 1274.020 0.090 1277.900 2.700 ;
        RECT 1279.620 0.090 1283.500 2.700 ;
        RECT 1285.220 0.090 1289.100 2.700 ;
        RECT 1290.820 0.090 1294.700 2.700 ;
        RECT 1296.420 0.090 1300.300 2.700 ;
        RECT 1302.020 0.090 1305.900 2.700 ;
        RECT 1307.620 0.090 1311.500 2.700 ;
        RECT 1313.220 0.090 1317.100 2.700 ;
        RECT 1318.820 0.090 1322.700 2.700 ;
        RECT 1324.420 0.090 1328.300 2.700 ;
        RECT 1330.020 0.090 1333.900 2.700 ;
        RECT 1335.620 0.090 1339.500 2.700 ;
        RECT 1341.220 0.090 1345.100 2.700 ;
        RECT 1346.820 0.090 1350.700 2.700 ;
        RECT 1352.420 0.090 1356.300 2.700 ;
        RECT 1358.020 0.090 1361.900 2.700 ;
        RECT 1363.620 0.090 1367.500 2.700 ;
        RECT 1369.220 0.090 1373.100 2.700 ;
        RECT 1374.820 0.090 1378.700 2.700 ;
        RECT 1380.420 0.090 1384.300 2.700 ;
        RECT 1386.020 0.090 1389.900 2.700 ;
        RECT 1391.620 0.090 1395.500 2.700 ;
        RECT 1397.220 0.090 1401.100 2.700 ;
        RECT 1402.820 0.090 1406.700 2.700 ;
        RECT 1408.420 0.090 1412.300 2.700 ;
        RECT 1414.020 0.090 1417.900 2.700 ;
        RECT 1419.620 0.090 1423.500 2.700 ;
        RECT 1425.220 0.090 1429.100 2.700 ;
        RECT 1430.820 0.090 1434.700 2.700 ;
        RECT 1436.420 0.090 1440.300 2.700 ;
        RECT 1442.020 0.090 1445.900 2.700 ;
        RECT 1447.620 0.090 1451.500 2.700 ;
        RECT 1453.220 0.090 1457.100 2.700 ;
        RECT 1458.820 0.090 1462.700 2.700 ;
        RECT 1464.420 0.090 1468.300 2.700 ;
        RECT 1470.020 0.090 1473.900 2.700 ;
        RECT 1475.620 0.090 1479.500 2.700 ;
        RECT 1481.220 0.090 1485.100 2.700 ;
        RECT 1486.820 0.090 1490.700 2.700 ;
        RECT 1492.420 0.090 1496.300 2.700 ;
        RECT 1498.020 0.090 1501.900 2.700 ;
        RECT 1503.620 0.090 1507.500 2.700 ;
        RECT 1509.220 0.090 1513.100 2.700 ;
        RECT 1514.820 0.090 1518.700 2.700 ;
        RECT 1520.420 0.090 1524.300 2.700 ;
        RECT 1526.020 0.090 1529.900 2.700 ;
        RECT 1531.620 0.090 1535.500 2.700 ;
        RECT 1537.220 0.090 1541.100 2.700 ;
        RECT 1542.820 0.090 1546.700 2.700 ;
        RECT 1548.420 0.090 1552.300 2.700 ;
        RECT 1554.020 0.090 1557.900 2.700 ;
        RECT 1559.620 0.090 1563.500 2.700 ;
        RECT 1565.220 0.090 1569.100 2.700 ;
        RECT 1570.820 0.090 1574.700 2.700 ;
        RECT 1576.420 0.090 1580.300 2.700 ;
        RECT 1582.020 0.090 1585.900 2.700 ;
        RECT 1587.620 0.090 1591.500 2.700 ;
        RECT 1593.220 0.090 1597.100 2.700 ;
        RECT 1598.820 0.090 1602.700 2.700 ;
        RECT 1604.420 0.090 1608.300 2.700 ;
        RECT 1610.020 0.090 1613.900 2.700 ;
        RECT 1615.620 0.090 1619.500 2.700 ;
        RECT 1621.220 0.090 1625.100 2.700 ;
        RECT 1626.820 0.090 1630.700 2.700 ;
        RECT 1632.420 0.090 1636.300 2.700 ;
        RECT 1638.020 0.090 1641.900 2.700 ;
        RECT 1643.620 0.090 1647.500 2.700 ;
        RECT 1649.220 0.090 1653.100 2.700 ;
        RECT 1654.820 0.090 1658.700 2.700 ;
        RECT 1660.420 0.090 1664.300 2.700 ;
        RECT 1666.020 0.090 1669.900 2.700 ;
        RECT 1671.620 0.090 1675.500 2.700 ;
        RECT 1677.220 0.090 1681.100 2.700 ;
        RECT 1682.820 0.090 1686.700 2.700 ;
        RECT 1688.420 0.090 1692.300 2.700 ;
        RECT 1694.020 0.090 1697.900 2.700 ;
        RECT 1699.620 0.090 1703.500 2.700 ;
        RECT 1705.220 0.090 1709.100 2.700 ;
        RECT 1710.820 0.090 1714.700 2.700 ;
        RECT 1716.420 0.090 1720.300 2.700 ;
        RECT 1722.020 0.090 1725.900 2.700 ;
        RECT 1727.620 0.090 1731.500 2.700 ;
        RECT 1733.220 0.090 1737.100 2.700 ;
        RECT 1738.820 0.090 1742.700 2.700 ;
        RECT 1744.420 0.090 1748.300 2.700 ;
        RECT 1750.020 0.090 1753.900 2.700 ;
        RECT 1755.620 0.090 1759.500 2.700 ;
        RECT 1761.220 0.090 1765.100 2.700 ;
        RECT 1766.820 0.090 1770.700 2.700 ;
        RECT 1772.420 0.090 1776.300 2.700 ;
        RECT 1778.020 0.090 1781.900 2.700 ;
        RECT 1783.620 0.090 1787.500 2.700 ;
        RECT 1789.220 0.090 1793.100 2.700 ;
        RECT 1794.820 0.090 1798.700 2.700 ;
        RECT 1800.420 0.090 1804.300 2.700 ;
        RECT 1806.020 0.090 1809.900 2.700 ;
        RECT 1811.620 0.090 1815.500 2.700 ;
        RECT 1817.220 0.090 1821.100 2.700 ;
        RECT 1822.820 0.090 1826.700 2.700 ;
        RECT 1828.420 0.090 1832.300 2.700 ;
        RECT 1834.020 0.090 1837.900 2.700 ;
        RECT 1839.620 0.090 1843.500 2.700 ;
        RECT 1845.220 0.090 1849.100 2.700 ;
        RECT 1850.820 0.090 1854.700 2.700 ;
        RECT 1856.420 0.090 1860.300 2.700 ;
        RECT 1862.020 0.090 1865.900 2.700 ;
        RECT 1867.620 0.090 1871.500 2.700 ;
        RECT 1873.220 0.090 1877.100 2.700 ;
        RECT 1878.820 0.090 1882.700 2.700 ;
        RECT 1884.420 0.090 1888.300 2.700 ;
        RECT 1890.020 0.090 1893.900 2.700 ;
        RECT 1895.620 0.090 1899.500 2.700 ;
        RECT 1901.220 0.090 1905.100 2.700 ;
        RECT 1906.820 0.090 1910.700 2.700 ;
        RECT 1912.420 0.090 1916.300 2.700 ;
        RECT 1918.020 0.090 1921.900 2.700 ;
        RECT 1923.620 0.090 1927.500 2.700 ;
        RECT 1929.220 0.090 1933.100 2.700 ;
        RECT 1934.820 0.090 1938.700 2.700 ;
        RECT 1940.420 0.090 1944.300 2.700 ;
        RECT 1946.020 0.090 1949.900 2.700 ;
        RECT 1951.620 0.090 1955.500 2.700 ;
        RECT 1957.220 0.090 1961.100 2.700 ;
        RECT 1962.820 0.090 1966.700 2.700 ;
        RECT 1968.420 0.090 1972.300 2.700 ;
        RECT 1974.020 0.090 1977.900 2.700 ;
        RECT 1979.620 0.090 1983.500 2.700 ;
        RECT 1985.220 0.090 1989.100 2.700 ;
        RECT 1990.820 0.090 1994.700 2.700 ;
        RECT 1996.420 0.090 2000.300 2.700 ;
        RECT 2002.020 0.090 2005.900 2.700 ;
        RECT 2007.620 0.090 2011.500 2.700 ;
        RECT 2013.220 0.090 2017.100 2.700 ;
        RECT 2018.820 0.090 2022.700 2.700 ;
        RECT 2024.420 0.090 2028.300 2.700 ;
        RECT 2030.020 0.090 2033.900 2.700 ;
        RECT 2035.620 0.090 2039.500 2.700 ;
        RECT 2041.220 0.090 2045.100 2.700 ;
        RECT 2046.820 0.090 2050.700 2.700 ;
        RECT 2052.420 0.090 2056.300 2.700 ;
        RECT 2058.020 0.090 2061.900 2.700 ;
        RECT 2063.620 0.090 2067.500 2.700 ;
        RECT 2069.220 0.090 2073.100 2.700 ;
        RECT 2074.820 0.090 2078.700 2.700 ;
        RECT 2080.420 0.090 2084.300 2.700 ;
        RECT 2086.020 0.090 2089.900 2.700 ;
        RECT 2091.620 0.090 2095.500 2.700 ;
        RECT 2097.220 0.090 2101.100 2.700 ;
        RECT 2102.820 0.090 2106.700 2.700 ;
        RECT 2108.420 0.090 2112.300 2.700 ;
        RECT 2114.020 0.090 2117.900 2.700 ;
        RECT 2119.620 0.090 2123.500 2.700 ;
        RECT 2125.220 0.090 2129.100 2.700 ;
        RECT 2130.820 0.090 2134.700 2.700 ;
        RECT 2136.420 0.090 2140.300 2.700 ;
        RECT 2142.020 0.090 2145.900 2.700 ;
        RECT 2147.620 0.090 2151.500 2.700 ;
        RECT 2153.220 0.090 2157.100 2.700 ;
        RECT 2158.820 0.090 2162.700 2.700 ;
        RECT 2164.420 0.090 2168.300 2.700 ;
        RECT 2170.020 0.090 2173.900 2.700 ;
        RECT 2175.620 0.090 2179.500 2.700 ;
        RECT 2181.220 0.090 2185.100 2.700 ;
        RECT 2186.820 0.090 2190.700 2.700 ;
        RECT 2192.420 0.090 2196.300 2.700 ;
        RECT 2198.020 0.090 2201.900 2.700 ;
        RECT 2203.620 0.090 2207.500 2.700 ;
        RECT 2209.220 0.090 2213.100 2.700 ;
        RECT 2214.820 0.090 2218.700 2.700 ;
        RECT 2220.420 0.090 2224.300 2.700 ;
        RECT 2226.020 0.090 2229.900 2.700 ;
        RECT 2231.620 0.090 2235.500 2.700 ;
        RECT 2237.220 0.090 2241.100 2.700 ;
        RECT 2242.820 0.090 2246.700 2.700 ;
        RECT 2248.420 0.090 2252.300 2.700 ;
        RECT 2254.020 0.090 2257.900 2.700 ;
        RECT 2259.620 0.090 2263.500 2.700 ;
        RECT 2265.220 0.090 2269.100 2.700 ;
        RECT 2270.820 0.090 2274.700 2.700 ;
        RECT 2276.420 0.090 2280.300 2.700 ;
        RECT 2282.020 0.090 2285.900 2.700 ;
        RECT 2287.620 0.090 2291.500 2.700 ;
        RECT 2293.220 0.090 2297.100 2.700 ;
        RECT 2298.820 0.090 2302.700 2.700 ;
        RECT 2304.420 0.090 2308.300 2.700 ;
        RECT 2310.020 0.090 2313.900 2.700 ;
        RECT 2315.620 0.090 2319.500 2.700 ;
        RECT 2321.220 0.090 2325.100 2.700 ;
        RECT 2326.820 0.090 2330.700 2.700 ;
        RECT 2332.420 0.090 2336.300 2.700 ;
        RECT 2338.020 0.090 2341.900 2.700 ;
        RECT 2343.620 0.090 2347.500 2.700 ;
        RECT 2349.220 0.090 2353.100 2.700 ;
        RECT 2354.820 0.090 2358.700 2.700 ;
        RECT 2360.420 0.090 2364.300 2.700 ;
        RECT 2366.020 0.090 2369.900 2.700 ;
        RECT 2371.620 0.090 2375.500 2.700 ;
        RECT 2377.220 0.090 2381.100 2.700 ;
        RECT 2382.820 0.090 2386.700 2.700 ;
        RECT 2388.420 0.090 2392.300 2.700 ;
        RECT 2394.020 0.090 2397.900 2.700 ;
        RECT 2399.620 0.090 2403.500 2.700 ;
        RECT 2405.220 0.090 2409.100 2.700 ;
        RECT 2410.820 0.090 2414.700 2.700 ;
        RECT 2416.420 0.090 2420.300 2.700 ;
        RECT 2422.020 0.090 2425.900 2.700 ;
        RECT 2427.620 0.090 2431.500 2.700 ;
        RECT 2433.220 0.090 2437.100 2.700 ;
        RECT 2438.820 0.090 2442.700 2.700 ;
        RECT 2444.420 0.090 2448.300 2.700 ;
        RECT 2450.020 0.090 2453.900 2.700 ;
        RECT 2455.620 0.090 2459.500 2.700 ;
        RECT 2461.220 0.090 2465.100 2.700 ;
        RECT 2466.820 0.090 2470.700 2.700 ;
        RECT 2472.420 0.090 2476.300 2.700 ;
        RECT 2478.020 0.090 2481.900 2.700 ;
        RECT 2483.620 0.090 2487.500 2.700 ;
        RECT 2489.220 0.090 2493.100 2.700 ;
        RECT 2494.820 0.090 2498.700 2.700 ;
        RECT 2500.420 0.090 2504.300 2.700 ;
        RECT 2506.020 0.090 2509.900 2.700 ;
        RECT 2511.620 0.090 2515.500 2.700 ;
        RECT 2517.220 0.090 2521.100 2.700 ;
        RECT 2522.820 0.090 2526.700 2.700 ;
        RECT 2528.420 0.090 2532.300 2.700 ;
        RECT 2534.020 0.090 2537.900 2.700 ;
        RECT 2539.620 0.090 2543.500 2.700 ;
        RECT 2545.220 0.090 2549.100 2.700 ;
        RECT 2550.820 0.090 2554.700 2.700 ;
        RECT 2556.420 0.090 2560.300 2.700 ;
        RECT 2562.020 0.090 2565.900 2.700 ;
        RECT 2567.620 0.090 2571.500 2.700 ;
        RECT 2573.220 0.090 2577.100 2.700 ;
        RECT 2578.820 0.090 2582.700 2.700 ;
        RECT 2584.420 0.090 2588.300 2.700 ;
        RECT 2590.020 0.090 2593.900 2.700 ;
        RECT 2595.620 0.090 2599.500 2.700 ;
        RECT 2601.220 0.090 2605.100 2.700 ;
        RECT 2606.820 0.090 2610.700 2.700 ;
        RECT 2612.420 0.090 2616.300 2.700 ;
        RECT 2618.020 0.090 2621.900 2.700 ;
        RECT 2623.620 0.090 2627.500 2.700 ;
        RECT 2629.220 0.090 2633.100 2.700 ;
        RECT 2634.820 0.090 2638.700 2.700 ;
        RECT 2640.420 0.090 2644.300 2.700 ;
        RECT 2646.020 0.090 2649.900 2.700 ;
        RECT 2651.620 0.090 2655.500 2.700 ;
        RECT 2657.220 0.090 2661.100 2.700 ;
        RECT 2662.820 0.090 2666.700 2.700 ;
        RECT 2668.420 0.090 2672.300 2.700 ;
        RECT 2674.020 0.090 2677.900 2.700 ;
        RECT 2679.620 0.090 2683.500 2.700 ;
        RECT 2685.220 0.090 2689.100 2.700 ;
        RECT 2690.820 0.090 2694.700 2.700 ;
        RECT 2696.420 0.090 2700.300 2.700 ;
        RECT 2702.020 0.090 2705.900 2.700 ;
        RECT 2707.620 0.090 2711.500 2.700 ;
        RECT 2713.220 0.090 2717.100 2.700 ;
        RECT 2718.820 0.090 2722.700 2.700 ;
        RECT 2724.420 0.090 2728.300 2.700 ;
        RECT 2730.020 0.090 2733.900 2.700 ;
        RECT 2735.620 0.090 2739.500 2.700 ;
        RECT 2741.220 0.090 2745.100 2.700 ;
        RECT 2746.820 0.090 2750.700 2.700 ;
        RECT 2752.420 0.090 2756.300 2.700 ;
        RECT 2758.020 0.090 2761.900 2.700 ;
        RECT 2763.620 0.090 2767.500 2.700 ;
        RECT 2769.220 0.090 2773.100 2.700 ;
        RECT 2774.820 0.090 2778.700 2.700 ;
        RECT 2780.420 0.090 2784.300 2.700 ;
        RECT 2786.020 0.090 2789.900 2.700 ;
        RECT 2791.620 0.090 2795.500 2.700 ;
        RECT 2797.220 0.090 2801.100 2.700 ;
        RECT 2802.820 0.090 2806.700 2.700 ;
        RECT 2808.420 0.090 2812.300 2.700 ;
        RECT 2814.020 0.090 2817.900 2.700 ;
        RECT 2819.620 0.090 2823.500 2.700 ;
        RECT 2825.220 0.090 2829.100 2.700 ;
        RECT 2830.820 0.090 2834.700 2.700 ;
        RECT 2836.420 0.090 2840.300 2.700 ;
        RECT 2842.020 0.090 2845.900 2.700 ;
        RECT 2847.620 0.090 2851.500 2.700 ;
        RECT 2853.220 0.090 2857.100 2.700 ;
        RECT 2858.820 0.090 2862.700 2.700 ;
        RECT 2864.420 0.090 2868.300 2.700 ;
        RECT 2870.020 0.090 2873.900 2.700 ;
        RECT 2875.620 0.090 2879.500 2.700 ;
        RECT 2881.220 0.090 2980.740 2.700 ;
      LAYER Metal3 ;
        RECT 1.820 2971.380 2998.100 2991.380 ;
        RECT 1.820 2969.700 2997.300 2971.380 ;
        RECT 2.700 2969.660 2997.300 2969.700 ;
        RECT 2.700 2967.980 2998.100 2969.660 ;
        RECT 1.820 2914.820 2998.100 2967.980 ;
        RECT 1.820 2914.260 2997.300 2914.820 ;
        RECT 2.700 2913.100 2997.300 2914.260 ;
        RECT 2.700 2912.540 2998.100 2913.100 ;
        RECT 1.820 2858.820 2998.100 2912.540 ;
        RECT 2.700 2858.260 2998.100 2858.820 ;
        RECT 2.700 2857.100 2997.300 2858.260 ;
        RECT 1.820 2856.540 2997.300 2857.100 ;
        RECT 1.820 2803.380 2998.100 2856.540 ;
        RECT 2.700 2801.700 2998.100 2803.380 ;
        RECT 2.700 2801.660 2997.300 2801.700 ;
        RECT 1.820 2799.980 2997.300 2801.660 ;
        RECT 1.820 2747.940 2998.100 2799.980 ;
        RECT 2.700 2746.220 2998.100 2747.940 ;
        RECT 1.820 2745.140 2998.100 2746.220 ;
        RECT 1.820 2743.420 2997.300 2745.140 ;
        RECT 1.820 2692.500 2998.100 2743.420 ;
        RECT 2.700 2690.780 2998.100 2692.500 ;
        RECT 1.820 2688.580 2998.100 2690.780 ;
        RECT 1.820 2686.860 2997.300 2688.580 ;
        RECT 1.820 2637.060 2998.100 2686.860 ;
        RECT 2.700 2635.340 2998.100 2637.060 ;
        RECT 1.820 2632.020 2998.100 2635.340 ;
        RECT 1.820 2630.300 2997.300 2632.020 ;
        RECT 1.820 2581.620 2998.100 2630.300 ;
        RECT 2.700 2579.900 2998.100 2581.620 ;
        RECT 1.820 2575.460 2998.100 2579.900 ;
        RECT 1.820 2573.740 2997.300 2575.460 ;
        RECT 1.820 2526.180 2998.100 2573.740 ;
        RECT 2.700 2524.460 2998.100 2526.180 ;
        RECT 1.820 2518.900 2998.100 2524.460 ;
        RECT 1.820 2517.180 2997.300 2518.900 ;
        RECT 1.820 2470.740 2998.100 2517.180 ;
        RECT 2.700 2469.020 2998.100 2470.740 ;
        RECT 1.820 2462.340 2998.100 2469.020 ;
        RECT 1.820 2460.620 2997.300 2462.340 ;
        RECT 1.820 2415.300 2998.100 2460.620 ;
        RECT 2.700 2413.580 2998.100 2415.300 ;
        RECT 1.820 2405.780 2998.100 2413.580 ;
        RECT 1.820 2404.060 2997.300 2405.780 ;
        RECT 1.820 2359.860 2998.100 2404.060 ;
        RECT 2.700 2358.140 2998.100 2359.860 ;
        RECT 1.820 2349.220 2998.100 2358.140 ;
        RECT 1.820 2347.500 2997.300 2349.220 ;
        RECT 1.820 2304.420 2998.100 2347.500 ;
        RECT 2.700 2302.700 2998.100 2304.420 ;
        RECT 1.820 2292.660 2998.100 2302.700 ;
        RECT 1.820 2290.940 2997.300 2292.660 ;
        RECT 1.820 2248.980 2998.100 2290.940 ;
        RECT 2.700 2247.260 2998.100 2248.980 ;
        RECT 1.820 2236.100 2998.100 2247.260 ;
        RECT 1.820 2234.380 2997.300 2236.100 ;
        RECT 1.820 2193.540 2998.100 2234.380 ;
        RECT 2.700 2191.820 2998.100 2193.540 ;
        RECT 1.820 2179.540 2998.100 2191.820 ;
        RECT 1.820 2177.820 2997.300 2179.540 ;
        RECT 1.820 2138.100 2998.100 2177.820 ;
        RECT 2.700 2136.380 2998.100 2138.100 ;
        RECT 1.820 2122.980 2998.100 2136.380 ;
        RECT 1.820 2121.260 2997.300 2122.980 ;
        RECT 1.820 2082.660 2998.100 2121.260 ;
        RECT 2.700 2080.940 2998.100 2082.660 ;
        RECT 1.820 2066.420 2998.100 2080.940 ;
        RECT 1.820 2064.700 2997.300 2066.420 ;
        RECT 1.820 2027.220 2998.100 2064.700 ;
        RECT 2.700 2025.500 2998.100 2027.220 ;
        RECT 1.820 2009.860 2998.100 2025.500 ;
        RECT 1.820 2008.140 2997.300 2009.860 ;
        RECT 1.820 1971.780 2998.100 2008.140 ;
        RECT 2.700 1970.060 2998.100 1971.780 ;
        RECT 1.820 1953.300 2998.100 1970.060 ;
        RECT 1.820 1951.580 2997.300 1953.300 ;
        RECT 1.820 1916.340 2998.100 1951.580 ;
        RECT 2.700 1914.620 2998.100 1916.340 ;
        RECT 1.820 1896.740 2998.100 1914.620 ;
        RECT 1.820 1895.020 2997.300 1896.740 ;
        RECT 1.820 1860.900 2998.100 1895.020 ;
        RECT 2.700 1859.180 2998.100 1860.900 ;
        RECT 1.820 1840.180 2998.100 1859.180 ;
        RECT 1.820 1838.460 2997.300 1840.180 ;
        RECT 1.820 1805.460 2998.100 1838.460 ;
        RECT 2.700 1803.740 2998.100 1805.460 ;
        RECT 1.820 1783.620 2998.100 1803.740 ;
        RECT 1.820 1781.900 2997.300 1783.620 ;
        RECT 1.820 1750.020 2998.100 1781.900 ;
        RECT 2.700 1748.300 2998.100 1750.020 ;
        RECT 1.820 1727.060 2998.100 1748.300 ;
        RECT 1.820 1725.340 2997.300 1727.060 ;
        RECT 1.820 1694.580 2998.100 1725.340 ;
        RECT 2.700 1692.860 2998.100 1694.580 ;
        RECT 1.820 1670.500 2998.100 1692.860 ;
        RECT 1.820 1668.780 2997.300 1670.500 ;
        RECT 1.820 1639.140 2998.100 1668.780 ;
        RECT 2.700 1637.420 2998.100 1639.140 ;
        RECT 1.820 1613.940 2998.100 1637.420 ;
        RECT 1.820 1612.220 2997.300 1613.940 ;
        RECT 1.820 1583.700 2998.100 1612.220 ;
        RECT 2.700 1581.980 2998.100 1583.700 ;
        RECT 1.820 1557.380 2998.100 1581.980 ;
        RECT 1.820 1555.660 2997.300 1557.380 ;
        RECT 1.820 1528.260 2998.100 1555.660 ;
        RECT 2.700 1526.540 2998.100 1528.260 ;
        RECT 1.820 1500.820 2998.100 1526.540 ;
        RECT 1.820 1499.100 2997.300 1500.820 ;
        RECT 1.820 1472.820 2998.100 1499.100 ;
        RECT 2.700 1471.100 2998.100 1472.820 ;
        RECT 1.820 1444.260 2998.100 1471.100 ;
        RECT 1.820 1442.540 2997.300 1444.260 ;
        RECT 1.820 1417.380 2998.100 1442.540 ;
        RECT 2.700 1415.660 2998.100 1417.380 ;
        RECT 1.820 1387.700 2998.100 1415.660 ;
        RECT 1.820 1385.980 2997.300 1387.700 ;
        RECT 1.820 1361.940 2998.100 1385.980 ;
        RECT 2.700 1360.220 2998.100 1361.940 ;
        RECT 1.820 1331.140 2998.100 1360.220 ;
        RECT 1.820 1329.420 2997.300 1331.140 ;
        RECT 1.820 1306.500 2998.100 1329.420 ;
        RECT 2.700 1304.780 2998.100 1306.500 ;
        RECT 1.820 1274.580 2998.100 1304.780 ;
        RECT 1.820 1272.860 2997.300 1274.580 ;
        RECT 1.820 1251.060 2998.100 1272.860 ;
        RECT 2.700 1249.340 2998.100 1251.060 ;
        RECT 1.820 1218.020 2998.100 1249.340 ;
        RECT 1.820 1216.300 2997.300 1218.020 ;
        RECT 1.820 1195.620 2998.100 1216.300 ;
        RECT 2.700 1193.900 2998.100 1195.620 ;
        RECT 1.820 1161.460 2998.100 1193.900 ;
        RECT 1.820 1159.740 2997.300 1161.460 ;
        RECT 1.820 1140.180 2998.100 1159.740 ;
        RECT 2.700 1138.460 2998.100 1140.180 ;
        RECT 1.820 1104.900 2998.100 1138.460 ;
        RECT 1.820 1103.180 2997.300 1104.900 ;
        RECT 1.820 1084.740 2998.100 1103.180 ;
        RECT 2.700 1083.020 2998.100 1084.740 ;
        RECT 1.820 1048.340 2998.100 1083.020 ;
        RECT 1.820 1046.620 2997.300 1048.340 ;
        RECT 1.820 1029.300 2998.100 1046.620 ;
        RECT 2.700 1027.580 2998.100 1029.300 ;
        RECT 1.820 991.780 2998.100 1027.580 ;
        RECT 1.820 990.060 2997.300 991.780 ;
        RECT 1.820 973.860 2998.100 990.060 ;
        RECT 2.700 972.140 2998.100 973.860 ;
        RECT 1.820 935.220 2998.100 972.140 ;
        RECT 1.820 933.500 2997.300 935.220 ;
        RECT 1.820 918.420 2998.100 933.500 ;
        RECT 2.700 916.700 2998.100 918.420 ;
        RECT 1.820 878.660 2998.100 916.700 ;
        RECT 1.820 876.940 2997.300 878.660 ;
        RECT 1.820 862.980 2998.100 876.940 ;
        RECT 2.700 861.260 2998.100 862.980 ;
        RECT 1.820 822.100 2998.100 861.260 ;
        RECT 1.820 820.380 2997.300 822.100 ;
        RECT 1.820 807.540 2998.100 820.380 ;
        RECT 2.700 805.820 2998.100 807.540 ;
        RECT 1.820 765.540 2998.100 805.820 ;
        RECT 1.820 763.820 2997.300 765.540 ;
        RECT 1.820 752.100 2998.100 763.820 ;
        RECT 2.700 750.380 2998.100 752.100 ;
        RECT 1.820 708.980 2998.100 750.380 ;
        RECT 1.820 707.260 2997.300 708.980 ;
        RECT 1.820 696.660 2998.100 707.260 ;
        RECT 2.700 694.940 2998.100 696.660 ;
        RECT 1.820 652.420 2998.100 694.940 ;
        RECT 1.820 650.700 2997.300 652.420 ;
        RECT 1.820 641.220 2998.100 650.700 ;
        RECT 2.700 639.500 2998.100 641.220 ;
        RECT 1.820 595.860 2998.100 639.500 ;
        RECT 1.820 594.140 2997.300 595.860 ;
        RECT 1.820 585.780 2998.100 594.140 ;
        RECT 2.700 584.060 2998.100 585.780 ;
        RECT 1.820 539.300 2998.100 584.060 ;
        RECT 1.820 537.580 2997.300 539.300 ;
        RECT 1.820 530.340 2998.100 537.580 ;
        RECT 2.700 528.620 2998.100 530.340 ;
        RECT 1.820 482.740 2998.100 528.620 ;
        RECT 1.820 481.020 2997.300 482.740 ;
        RECT 1.820 474.900 2998.100 481.020 ;
        RECT 2.700 473.180 2998.100 474.900 ;
        RECT 1.820 426.180 2998.100 473.180 ;
        RECT 1.820 424.460 2997.300 426.180 ;
        RECT 1.820 419.460 2998.100 424.460 ;
        RECT 2.700 417.740 2998.100 419.460 ;
        RECT 1.820 369.620 2998.100 417.740 ;
        RECT 1.820 367.900 2997.300 369.620 ;
        RECT 1.820 364.020 2998.100 367.900 ;
        RECT 2.700 362.300 2998.100 364.020 ;
        RECT 1.820 313.060 2998.100 362.300 ;
        RECT 1.820 311.340 2997.300 313.060 ;
        RECT 1.820 308.580 2998.100 311.340 ;
        RECT 2.700 306.860 2998.100 308.580 ;
        RECT 1.820 256.500 2998.100 306.860 ;
        RECT 1.820 254.780 2997.300 256.500 ;
        RECT 1.820 253.140 2998.100 254.780 ;
        RECT 2.700 251.420 2998.100 253.140 ;
        RECT 1.820 199.940 2998.100 251.420 ;
        RECT 1.820 198.220 2997.300 199.940 ;
        RECT 1.820 197.700 2998.100 198.220 ;
        RECT 2.700 195.980 2998.100 197.700 ;
        RECT 1.820 143.380 2998.100 195.980 ;
        RECT 1.820 142.260 2997.300 143.380 ;
        RECT 2.700 141.660 2997.300 142.260 ;
        RECT 2.700 140.540 2998.100 141.660 ;
        RECT 1.820 86.820 2998.100 140.540 ;
        RECT 2.700 85.100 2997.300 86.820 ;
        RECT 1.820 31.380 2998.100 85.100 ;
        RECT 2.700 30.260 2998.100 31.380 ;
        RECT 2.700 29.660 2997.300 30.260 ;
        RECT 1.820 28.540 2997.300 29.660 ;
        RECT 1.820 0.140 2998.100 28.540 ;
      LAYER Metal4 ;
        RECT 609.370 2334.970 624.270 2341.830 ;
        RECT 627.970 2334.970 642.870 2341.830 ;
        RECT 646.570 2334.970 661.470 2341.830 ;
        RECT 665.170 2334.970 680.070 2341.830 ;
        RECT 683.770 2334.970 729.870 2341.830 ;
        RECT 733.570 2334.970 748.470 2341.830 ;
        RECT 752.170 2334.970 767.070 2341.830 ;
        RECT 770.770 2334.970 785.670 2341.830 ;
        RECT 789.370 2334.970 804.270 2341.830 ;
        RECT 807.970 2334.970 822.870 2341.830 ;
        RECT 826.570 2337.040 841.470 2341.830 ;
        RECT 845.170 2337.040 860.070 2341.830 ;
        RECT 826.570 2334.970 860.070 2337.040 ;
        RECT 863.770 2334.970 909.870 2341.830 ;
        RECT 913.570 2334.970 928.470 2341.830 ;
        RECT 932.170 2334.970 947.070 2341.830 ;
        RECT 950.770 2334.970 965.670 2341.830 ;
        RECT 969.370 2334.970 984.270 2341.830 ;
        RECT 987.970 2334.970 1002.870 2341.830 ;
        RECT 1006.570 2334.970 1021.470 2341.830 ;
        RECT 1025.170 2334.970 1040.070 2341.830 ;
        RECT 1043.770 2334.970 1089.870 2341.830 ;
        RECT 1093.570 2334.970 1108.470 2341.830 ;
        RECT 1112.170 2334.970 1127.070 2341.830 ;
        RECT 1130.770 2337.040 1145.670 2341.830 ;
        RECT 1149.370 2337.040 1164.270 2341.830 ;
        RECT 1130.770 2334.970 1164.270 2337.040 ;
        RECT 1167.970 2334.970 1182.870 2341.830 ;
        RECT 1186.570 2334.970 1201.470 2341.830 ;
        RECT 1205.170 2334.970 1220.070 2341.830 ;
        RECT 1223.770 2334.970 1269.870 2341.830 ;
        RECT 1273.570 2334.970 1288.470 2341.830 ;
        RECT 1292.170 2334.970 1307.070 2341.830 ;
        RECT 1310.770 2334.970 1325.670 2341.830 ;
        RECT 1329.370 2334.970 1344.270 2341.830 ;
        RECT 1347.970 2334.970 1362.870 2341.830 ;
        RECT 1366.570 2334.970 1381.470 2341.830 ;
        RECT 1385.170 2334.970 1400.070 2341.830 ;
        RECT 1403.770 2334.970 1449.870 2341.830 ;
        RECT 1453.570 2334.970 1468.470 2341.830 ;
        RECT 1472.170 2334.970 1487.070 2341.830 ;
        RECT 1490.770 2334.970 1505.670 2341.830 ;
        RECT 1509.370 2334.970 1524.270 2341.830 ;
        RECT 1527.970 2334.970 1542.870 2341.830 ;
        RECT 1546.570 2334.970 1561.470 2341.830 ;
        RECT 1565.170 2334.970 1580.070 2341.830 ;
        RECT 1583.770 2334.970 1629.870 2341.830 ;
        RECT 1633.570 2334.970 1648.470 2341.830 ;
        RECT 1652.170 2334.970 1667.070 2341.830 ;
        RECT 1670.770 2337.040 1685.670 2341.830 ;
        RECT 1689.370 2337.040 1704.270 2341.830 ;
        RECT 1670.770 2334.970 1704.270 2337.040 ;
        RECT 1707.970 2334.970 1722.870 2341.830 ;
        RECT 1726.570 2334.970 1741.470 2341.830 ;
        RECT 1745.170 2337.040 1760.070 2341.830 ;
        RECT 1763.770 2337.040 1809.870 2341.830 ;
        RECT 1745.170 2334.970 1809.870 2337.040 ;
        RECT 1813.570 2334.970 1828.470 2341.830 ;
        RECT 1832.170 2334.970 1847.070 2341.830 ;
        RECT 1850.770 2334.970 1865.670 2341.830 ;
        RECT 1869.370 2334.970 1884.270 2341.830 ;
        RECT 1887.970 2334.970 1902.870 2341.830 ;
        RECT 1906.570 2334.970 1921.470 2341.830 ;
        RECT 1925.170 2334.970 1940.070 2341.830 ;
        RECT 1943.770 2337.040 1989.870 2341.830 ;
        RECT 1993.570 2337.040 2008.470 2341.830 ;
        RECT 1943.770 2334.970 2008.470 2337.040 ;
        RECT 2012.170 2334.970 2027.070 2341.830 ;
        RECT 608.360 851.380 2027.070 2334.970 ;
        RECT 608.360 851.350 661.470 851.380 ;
        RECT 609.370 20.250 624.270 851.350 ;
        RECT 627.970 20.250 642.870 851.350 ;
        RECT 646.570 20.250 661.470 851.350 ;
        RECT 665.170 851.350 1021.470 851.380 ;
        RECT 665.170 20.250 680.070 851.350 ;
        RECT 683.770 20.250 729.870 851.350 ;
        RECT 733.570 20.250 748.470 851.350 ;
        RECT 752.170 20.250 767.070 851.350 ;
        RECT 770.770 20.250 785.670 851.350 ;
        RECT 789.370 20.250 804.270 851.350 ;
        RECT 807.970 20.250 822.870 851.350 ;
        RECT 826.570 850.400 860.070 851.350 ;
        RECT 826.570 20.250 841.470 850.400 ;
        RECT 845.170 20.250 860.070 850.400 ;
        RECT 863.770 20.250 909.870 851.350 ;
        RECT 913.570 20.250 928.470 851.350 ;
        RECT 932.170 20.250 947.070 851.350 ;
        RECT 950.770 20.250 965.670 851.350 ;
        RECT 969.370 20.250 984.270 851.350 ;
        RECT 987.970 20.250 1002.870 851.350 ;
        RECT 1006.570 20.250 1021.470 851.350 ;
        RECT 1025.170 851.350 1201.470 851.380 ;
        RECT 1025.170 20.250 1040.070 851.350 ;
        RECT 1043.770 20.250 1089.870 851.350 ;
        RECT 1093.570 20.250 1108.470 851.350 ;
        RECT 1112.170 20.250 1127.070 851.350 ;
        RECT 1130.770 850.400 1164.270 851.350 ;
        RECT 1130.770 20.250 1145.670 850.400 ;
        RECT 1149.370 20.250 1164.270 850.400 ;
        RECT 1167.970 20.250 1182.870 851.350 ;
        RECT 1186.570 20.250 1201.470 851.350 ;
        RECT 1205.170 851.350 1381.470 851.380 ;
        RECT 1205.170 20.250 1220.070 851.350 ;
        RECT 1223.770 20.250 1269.870 851.350 ;
        RECT 1273.570 20.250 1288.470 851.350 ;
        RECT 1292.170 20.250 1307.070 851.350 ;
        RECT 1310.770 20.250 1325.670 851.350 ;
        RECT 1329.370 20.250 1344.270 851.350 ;
        RECT 1347.970 20.250 1362.870 851.350 ;
        RECT 1366.570 20.250 1381.470 851.350 ;
        RECT 1385.170 851.350 1561.470 851.380 ;
        RECT 1385.170 20.250 1400.070 851.350 ;
        RECT 1403.770 20.250 1449.870 851.350 ;
        RECT 1453.570 20.250 1468.470 851.350 ;
        RECT 1472.170 20.250 1487.070 851.350 ;
        RECT 1490.770 20.250 1505.670 851.350 ;
        RECT 1509.370 20.250 1524.270 851.350 ;
        RECT 1527.970 20.250 1542.870 851.350 ;
        RECT 1546.570 20.250 1561.470 851.350 ;
        RECT 1565.170 851.350 1741.470 851.380 ;
        RECT 1565.170 20.250 1580.070 851.350 ;
        RECT 1583.770 20.250 1629.870 851.350 ;
        RECT 1633.570 20.250 1648.470 851.350 ;
        RECT 1652.170 20.250 1667.070 851.350 ;
        RECT 1670.770 850.400 1704.270 851.350 ;
        RECT 1670.770 20.250 1685.670 850.400 ;
        RECT 1689.370 20.250 1704.270 850.400 ;
        RECT 1707.970 20.250 1722.870 851.350 ;
        RECT 1726.570 20.250 1741.470 851.350 ;
        RECT 1745.170 851.350 1921.470 851.380 ;
        RECT 1745.170 850.400 1809.870 851.350 ;
        RECT 1745.170 20.250 1760.070 850.400 ;
        RECT 1763.770 20.250 1809.870 850.400 ;
        RECT 1813.570 20.250 1828.470 851.350 ;
        RECT 1832.170 20.250 1847.070 851.350 ;
        RECT 1850.770 20.250 1865.670 851.350 ;
        RECT 1869.370 20.250 1884.270 851.350 ;
        RECT 1887.970 20.250 1902.870 851.350 ;
        RECT 1906.570 20.250 1921.470 851.350 ;
        RECT 1925.170 851.350 2027.070 851.380 ;
        RECT 1925.170 20.250 1940.070 851.350 ;
        RECT 1943.770 850.400 2008.470 851.350 ;
        RECT 1943.770 20.250 1989.870 850.400 ;
        RECT 1993.570 20.250 2008.470 850.400 ;
        RECT 2012.170 20.250 2027.070 851.350 ;
        RECT 2030.770 20.250 2045.670 2341.830 ;
        RECT 2049.370 20.250 2064.270 2341.830 ;
        RECT 2067.970 20.250 2070.540 2341.830 ;
      LAYER Metal5 ;
        RECT 608.280 1019.220 1986.320 2285.260 ;
  END
END user_project_wrapper
END LIBRARY

